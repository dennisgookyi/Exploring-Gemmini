module cc_dir_ext(
  input  [9:0]   RW0_addr,
  input          RW0_clk,
  input  [135:0] RW0_wdata,
  output [135:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [7:0]   RW0_wmask
);
  wire [9:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [16:0] mem_0_0_RW0_wdata;
  wire [16:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [9:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [16:0] mem_0_1_RW0_wdata;
  wire [16:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [9:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [16:0] mem_0_2_RW0_wdata;
  wire [16:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [9:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [16:0] mem_0_3_RW0_wdata;
  wire [16:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [9:0] mem_0_4_RW0_addr;
  wire  mem_0_4_RW0_clk;
  wire [16:0] mem_0_4_RW0_wdata;
  wire [16:0] mem_0_4_RW0_rdata;
  wire  mem_0_4_RW0_en;
  wire  mem_0_4_RW0_wmode;
  wire  mem_0_4_RW0_wmask;
  wire [9:0] mem_0_5_RW0_addr;
  wire  mem_0_5_RW0_clk;
  wire [16:0] mem_0_5_RW0_wdata;
  wire [16:0] mem_0_5_RW0_rdata;
  wire  mem_0_5_RW0_en;
  wire  mem_0_5_RW0_wmode;
  wire  mem_0_5_RW0_wmask;
  wire [9:0] mem_0_6_RW0_addr;
  wire  mem_0_6_RW0_clk;
  wire [16:0] mem_0_6_RW0_wdata;
  wire [16:0] mem_0_6_RW0_rdata;
  wire  mem_0_6_RW0_en;
  wire  mem_0_6_RW0_wmode;
  wire  mem_0_6_RW0_wmask;
  wire [9:0] mem_0_7_RW0_addr;
  wire  mem_0_7_RW0_clk;
  wire [16:0] mem_0_7_RW0_wdata;
  wire [16:0] mem_0_7_RW0_rdata;
  wire  mem_0_7_RW0_en;
  wire  mem_0_7_RW0_wmode;
  wire  mem_0_7_RW0_wmask;
  wire [16:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [16:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [16:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [16:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [16:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata;
  wire [16:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata;
  wire [16:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata;
  wire [16:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata;
  wire [33:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [50:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [67:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [84:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [101:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [118:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [135:0] RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [33:0] _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [50:0] _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [67:0] _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [84:0] _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [101:0] _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [118:0] _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  split_cc_dir_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 (
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 (
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 (
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 (
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[16:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[33:17];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[50:34];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[67:51];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_RW0_addr = RW0_addr;
  assign mem_0_4_RW0_clk = RW0_clk;
  assign mem_0_4_RW0_wdata = RW0_wdata[84:68];
  assign mem_0_4_RW0_en = RW0_en;
  assign mem_0_4_RW0_wmode = RW0_wmode;
  assign mem_0_4_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_RW0_addr = RW0_addr;
  assign mem_0_5_RW0_clk = RW0_clk;
  assign mem_0_5_RW0_wdata = RW0_wdata[101:85];
  assign mem_0_5_RW0_en = RW0_en;
  assign mem_0_5_RW0_wmode = RW0_wmode;
  assign mem_0_5_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_RW0_addr = RW0_addr;
  assign mem_0_6_RW0_clk = RW0_clk;
  assign mem_0_6_RW0_wdata = RW0_wdata[118:102];
  assign mem_0_6_RW0_en = RW0_en;
  assign mem_0_6_RW0_wmode = RW0_wmode;
  assign mem_0_6_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_RW0_addr = RW0_addr;
  assign mem_0_7_RW0_clk = RW0_clk;
  assign mem_0_7_RW0_wdata = RW0_wdata[135:119];
  assign mem_0_7_RW0_en = RW0_en;
  assign mem_0_7_RW0_wmode = RW0_wmode;
  assign mem_0_7_RW0_wmask = RW0_wmask[7];
endmodule
module cc_banks_0_ext(
  input  [12:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [12:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [63:0] mem_0_0_RW0_wdata;
  wire [63:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0;
  split_cc_banks_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata;
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata;
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
endmodule
module data_arrays_0_ext(
  input  [7:0]   RW0_addr,
  input          RW0_clk,
  input  [255:0] RW0_wdata,
  output [255:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [31:0]  RW0_wmask
);
  wire [7:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [7:0] mem_0_0_RW0_wdata;
  wire [7:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [7:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [7:0] mem_0_1_RW0_wdata;
  wire [7:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [7:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [7:0] mem_0_2_RW0_wdata;
  wire [7:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [7:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [7:0] mem_0_3_RW0_wdata;
  wire [7:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [7:0] mem_0_4_RW0_addr;
  wire  mem_0_4_RW0_clk;
  wire [7:0] mem_0_4_RW0_wdata;
  wire [7:0] mem_0_4_RW0_rdata;
  wire  mem_0_4_RW0_en;
  wire  mem_0_4_RW0_wmode;
  wire  mem_0_4_RW0_wmask;
  wire [7:0] mem_0_5_RW0_addr;
  wire  mem_0_5_RW0_clk;
  wire [7:0] mem_0_5_RW0_wdata;
  wire [7:0] mem_0_5_RW0_rdata;
  wire  mem_0_5_RW0_en;
  wire  mem_0_5_RW0_wmode;
  wire  mem_0_5_RW0_wmask;
  wire [7:0] mem_0_6_RW0_addr;
  wire  mem_0_6_RW0_clk;
  wire [7:0] mem_0_6_RW0_wdata;
  wire [7:0] mem_0_6_RW0_rdata;
  wire  mem_0_6_RW0_en;
  wire  mem_0_6_RW0_wmode;
  wire  mem_0_6_RW0_wmask;
  wire [7:0] mem_0_7_RW0_addr;
  wire  mem_0_7_RW0_clk;
  wire [7:0] mem_0_7_RW0_wdata;
  wire [7:0] mem_0_7_RW0_rdata;
  wire  mem_0_7_RW0_en;
  wire  mem_0_7_RW0_wmode;
  wire  mem_0_7_RW0_wmask;
  wire [7:0] mem_0_8_RW0_addr;
  wire  mem_0_8_RW0_clk;
  wire [7:0] mem_0_8_RW0_wdata;
  wire [7:0] mem_0_8_RW0_rdata;
  wire  mem_0_8_RW0_en;
  wire  mem_0_8_RW0_wmode;
  wire  mem_0_8_RW0_wmask;
  wire [7:0] mem_0_9_RW0_addr;
  wire  mem_0_9_RW0_clk;
  wire [7:0] mem_0_9_RW0_wdata;
  wire [7:0] mem_0_9_RW0_rdata;
  wire  mem_0_9_RW0_en;
  wire  mem_0_9_RW0_wmode;
  wire  mem_0_9_RW0_wmask;
  wire [7:0] mem_0_10_RW0_addr;
  wire  mem_0_10_RW0_clk;
  wire [7:0] mem_0_10_RW0_wdata;
  wire [7:0] mem_0_10_RW0_rdata;
  wire  mem_0_10_RW0_en;
  wire  mem_0_10_RW0_wmode;
  wire  mem_0_10_RW0_wmask;
  wire [7:0] mem_0_11_RW0_addr;
  wire  mem_0_11_RW0_clk;
  wire [7:0] mem_0_11_RW0_wdata;
  wire [7:0] mem_0_11_RW0_rdata;
  wire  mem_0_11_RW0_en;
  wire  mem_0_11_RW0_wmode;
  wire  mem_0_11_RW0_wmask;
  wire [7:0] mem_0_12_RW0_addr;
  wire  mem_0_12_RW0_clk;
  wire [7:0] mem_0_12_RW0_wdata;
  wire [7:0] mem_0_12_RW0_rdata;
  wire  mem_0_12_RW0_en;
  wire  mem_0_12_RW0_wmode;
  wire  mem_0_12_RW0_wmask;
  wire [7:0] mem_0_13_RW0_addr;
  wire  mem_0_13_RW0_clk;
  wire [7:0] mem_0_13_RW0_wdata;
  wire [7:0] mem_0_13_RW0_rdata;
  wire  mem_0_13_RW0_en;
  wire  mem_0_13_RW0_wmode;
  wire  mem_0_13_RW0_wmask;
  wire [7:0] mem_0_14_RW0_addr;
  wire  mem_0_14_RW0_clk;
  wire [7:0] mem_0_14_RW0_wdata;
  wire [7:0] mem_0_14_RW0_rdata;
  wire  mem_0_14_RW0_en;
  wire  mem_0_14_RW0_wmode;
  wire  mem_0_14_RW0_wmask;
  wire [7:0] mem_0_15_RW0_addr;
  wire  mem_0_15_RW0_clk;
  wire [7:0] mem_0_15_RW0_wdata;
  wire [7:0] mem_0_15_RW0_rdata;
  wire  mem_0_15_RW0_en;
  wire  mem_0_15_RW0_wmode;
  wire  mem_0_15_RW0_wmask;
  wire [7:0] mem_0_16_RW0_addr;
  wire  mem_0_16_RW0_clk;
  wire [7:0] mem_0_16_RW0_wdata;
  wire [7:0] mem_0_16_RW0_rdata;
  wire  mem_0_16_RW0_en;
  wire  mem_0_16_RW0_wmode;
  wire  mem_0_16_RW0_wmask;
  wire [7:0] mem_0_17_RW0_addr;
  wire  mem_0_17_RW0_clk;
  wire [7:0] mem_0_17_RW0_wdata;
  wire [7:0] mem_0_17_RW0_rdata;
  wire  mem_0_17_RW0_en;
  wire  mem_0_17_RW0_wmode;
  wire  mem_0_17_RW0_wmask;
  wire [7:0] mem_0_18_RW0_addr;
  wire  mem_0_18_RW0_clk;
  wire [7:0] mem_0_18_RW0_wdata;
  wire [7:0] mem_0_18_RW0_rdata;
  wire  mem_0_18_RW0_en;
  wire  mem_0_18_RW0_wmode;
  wire  mem_0_18_RW0_wmask;
  wire [7:0] mem_0_19_RW0_addr;
  wire  mem_0_19_RW0_clk;
  wire [7:0] mem_0_19_RW0_wdata;
  wire [7:0] mem_0_19_RW0_rdata;
  wire  mem_0_19_RW0_en;
  wire  mem_0_19_RW0_wmode;
  wire  mem_0_19_RW0_wmask;
  wire [7:0] mem_0_20_RW0_addr;
  wire  mem_0_20_RW0_clk;
  wire [7:0] mem_0_20_RW0_wdata;
  wire [7:0] mem_0_20_RW0_rdata;
  wire  mem_0_20_RW0_en;
  wire  mem_0_20_RW0_wmode;
  wire  mem_0_20_RW0_wmask;
  wire [7:0] mem_0_21_RW0_addr;
  wire  mem_0_21_RW0_clk;
  wire [7:0] mem_0_21_RW0_wdata;
  wire [7:0] mem_0_21_RW0_rdata;
  wire  mem_0_21_RW0_en;
  wire  mem_0_21_RW0_wmode;
  wire  mem_0_21_RW0_wmask;
  wire [7:0] mem_0_22_RW0_addr;
  wire  mem_0_22_RW0_clk;
  wire [7:0] mem_0_22_RW0_wdata;
  wire [7:0] mem_0_22_RW0_rdata;
  wire  mem_0_22_RW0_en;
  wire  mem_0_22_RW0_wmode;
  wire  mem_0_22_RW0_wmask;
  wire [7:0] mem_0_23_RW0_addr;
  wire  mem_0_23_RW0_clk;
  wire [7:0] mem_0_23_RW0_wdata;
  wire [7:0] mem_0_23_RW0_rdata;
  wire  mem_0_23_RW0_en;
  wire  mem_0_23_RW0_wmode;
  wire  mem_0_23_RW0_wmask;
  wire [7:0] mem_0_24_RW0_addr;
  wire  mem_0_24_RW0_clk;
  wire [7:0] mem_0_24_RW0_wdata;
  wire [7:0] mem_0_24_RW0_rdata;
  wire  mem_0_24_RW0_en;
  wire  mem_0_24_RW0_wmode;
  wire  mem_0_24_RW0_wmask;
  wire [7:0] mem_0_25_RW0_addr;
  wire  mem_0_25_RW0_clk;
  wire [7:0] mem_0_25_RW0_wdata;
  wire [7:0] mem_0_25_RW0_rdata;
  wire  mem_0_25_RW0_en;
  wire  mem_0_25_RW0_wmode;
  wire  mem_0_25_RW0_wmask;
  wire [7:0] mem_0_26_RW0_addr;
  wire  mem_0_26_RW0_clk;
  wire [7:0] mem_0_26_RW0_wdata;
  wire [7:0] mem_0_26_RW0_rdata;
  wire  mem_0_26_RW0_en;
  wire  mem_0_26_RW0_wmode;
  wire  mem_0_26_RW0_wmask;
  wire [7:0] mem_0_27_RW0_addr;
  wire  mem_0_27_RW0_clk;
  wire [7:0] mem_0_27_RW0_wdata;
  wire [7:0] mem_0_27_RW0_rdata;
  wire  mem_0_27_RW0_en;
  wire  mem_0_27_RW0_wmode;
  wire  mem_0_27_RW0_wmask;
  wire [7:0] mem_0_28_RW0_addr;
  wire  mem_0_28_RW0_clk;
  wire [7:0] mem_0_28_RW0_wdata;
  wire [7:0] mem_0_28_RW0_rdata;
  wire  mem_0_28_RW0_en;
  wire  mem_0_28_RW0_wmode;
  wire  mem_0_28_RW0_wmask;
  wire [7:0] mem_0_29_RW0_addr;
  wire  mem_0_29_RW0_clk;
  wire [7:0] mem_0_29_RW0_wdata;
  wire [7:0] mem_0_29_RW0_rdata;
  wire  mem_0_29_RW0_en;
  wire  mem_0_29_RW0_wmode;
  wire  mem_0_29_RW0_wmask;
  wire [7:0] mem_0_30_RW0_addr;
  wire  mem_0_30_RW0_clk;
  wire [7:0] mem_0_30_RW0_wdata;
  wire [7:0] mem_0_30_RW0_rdata;
  wire  mem_0_30_RW0_en;
  wire  mem_0_30_RW0_wmode;
  wire  mem_0_30_RW0_wmask;
  wire [7:0] mem_0_31_RW0_addr;
  wire  mem_0_31_RW0_clk;
  wire [7:0] mem_0_31_RW0_wdata;
  wire [7:0] mem_0_31_RW0_rdata;
  wire  mem_0_31_RW0_en;
  wire  mem_0_31_RW0_wmode;
  wire  mem_0_31_RW0_wmask;
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [7:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata;
  wire [7:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata;
  wire [7:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata;
  wire [7:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata;
  wire [7:0] RW0_rdata_0_8 = mem_0_8_RW0_rdata;
  wire [7:0] RW0_rdata_0_9 = mem_0_9_RW0_rdata;
  wire [7:0] RW0_rdata_0_10 = mem_0_10_RW0_rdata;
  wire [7:0] RW0_rdata_0_11 = mem_0_11_RW0_rdata;
  wire [7:0] RW0_rdata_0_12 = mem_0_12_RW0_rdata;
  wire [7:0] RW0_rdata_0_13 = mem_0_13_RW0_rdata;
  wire [7:0] RW0_rdata_0_14 = mem_0_14_RW0_rdata;
  wire [7:0] RW0_rdata_0_15 = mem_0_15_RW0_rdata;
  wire [7:0] RW0_rdata_0_16 = mem_0_16_RW0_rdata;
  wire [7:0] RW0_rdata_0_17 = mem_0_17_RW0_rdata;
  wire [7:0] RW0_rdata_0_18 = mem_0_18_RW0_rdata;
  wire [7:0] RW0_rdata_0_19 = mem_0_19_RW0_rdata;
  wire [7:0] RW0_rdata_0_20 = mem_0_20_RW0_rdata;
  wire [7:0] RW0_rdata_0_21 = mem_0_21_RW0_rdata;
  wire [7:0] RW0_rdata_0_22 = mem_0_22_RW0_rdata;
  wire [7:0] RW0_rdata_0_23 = mem_0_23_RW0_rdata;
  wire [7:0] RW0_rdata_0_24 = mem_0_24_RW0_rdata;
  wire [7:0] RW0_rdata_0_25 = mem_0_25_RW0_rdata;
  wire [7:0] RW0_rdata_0_26 = mem_0_26_RW0_rdata;
  wire [7:0] RW0_rdata_0_27 = mem_0_27_RW0_rdata;
  wire [7:0] RW0_rdata_0_28 = mem_0_28_RW0_rdata;
  wire [7:0] RW0_rdata_0_29 = mem_0_29_RW0_rdata;
  wire [7:0] RW0_rdata_0_30 = mem_0_30_RW0_rdata;
  wire [7:0] RW0_rdata_0_31 = mem_0_31_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_6 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_7 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_8 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_9 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [127:0] _GEN_14 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8};
  wire [135:0] _GEN_15 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8};
  wire [143:0] _GEN_16 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [151:0] _GEN_17 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [159:0] _GEN_18 = {RW0_rdata_0_19,_GEN_17};
  wire [167:0] _GEN_19 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [175:0] _GEN_20 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [183:0] _GEN_21 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [191:0] _GEN_22 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [199:0] _GEN_23 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17};
  wire [207:0] _GEN_24 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17};
  wire [215:0] _GEN_25 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [223:0] _GEN_26 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [231:0] _GEN_27 = {RW0_rdata_0_28,_GEN_26};
  wire [239:0] _GEN_28 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [247:0] _GEN_29 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [255:0] RW0_rdata_0 = {RW0_rdata_0_31,RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [15:0] _GEN_30 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_31 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_32 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_33 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_34 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_35 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_36 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_37 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_38 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_39 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_40 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_41 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_42 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_43 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [127:0] _GEN_44 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8};
  wire [135:0] _GEN_45 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8};
  wire [143:0] _GEN_46 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [151:0] _GEN_47 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [159:0] _GEN_48 = {RW0_rdata_0_19,_GEN_17};
  wire [167:0] _GEN_49 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [175:0] _GEN_50 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [183:0] _GEN_51 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [191:0] _GEN_52 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [199:0] _GEN_53 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17};
  wire [207:0] _GEN_54 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17};
  wire [215:0] _GEN_55 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [223:0] _GEN_56 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [231:0] _GEN_57 = {RW0_rdata_0_28,_GEN_26};
  wire [239:0] _GEN_58 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [247:0] _GEN_59 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  split_data_arrays_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_4 (
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_5 (
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_6 (
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_7 (
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_8 (
    .RW0_addr(mem_0_8_RW0_addr),
    .RW0_clk(mem_0_8_RW0_clk),
    .RW0_wdata(mem_0_8_RW0_wdata),
    .RW0_rdata(mem_0_8_RW0_rdata),
    .RW0_en(mem_0_8_RW0_en),
    .RW0_wmode(mem_0_8_RW0_wmode),
    .RW0_wmask(mem_0_8_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_9 (
    .RW0_addr(mem_0_9_RW0_addr),
    .RW0_clk(mem_0_9_RW0_clk),
    .RW0_wdata(mem_0_9_RW0_wdata),
    .RW0_rdata(mem_0_9_RW0_rdata),
    .RW0_en(mem_0_9_RW0_en),
    .RW0_wmode(mem_0_9_RW0_wmode),
    .RW0_wmask(mem_0_9_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_10 (
    .RW0_addr(mem_0_10_RW0_addr),
    .RW0_clk(mem_0_10_RW0_clk),
    .RW0_wdata(mem_0_10_RW0_wdata),
    .RW0_rdata(mem_0_10_RW0_rdata),
    .RW0_en(mem_0_10_RW0_en),
    .RW0_wmode(mem_0_10_RW0_wmode),
    .RW0_wmask(mem_0_10_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_11 (
    .RW0_addr(mem_0_11_RW0_addr),
    .RW0_clk(mem_0_11_RW0_clk),
    .RW0_wdata(mem_0_11_RW0_wdata),
    .RW0_rdata(mem_0_11_RW0_rdata),
    .RW0_en(mem_0_11_RW0_en),
    .RW0_wmode(mem_0_11_RW0_wmode),
    .RW0_wmask(mem_0_11_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_12 (
    .RW0_addr(mem_0_12_RW0_addr),
    .RW0_clk(mem_0_12_RW0_clk),
    .RW0_wdata(mem_0_12_RW0_wdata),
    .RW0_rdata(mem_0_12_RW0_rdata),
    .RW0_en(mem_0_12_RW0_en),
    .RW0_wmode(mem_0_12_RW0_wmode),
    .RW0_wmask(mem_0_12_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_13 (
    .RW0_addr(mem_0_13_RW0_addr),
    .RW0_clk(mem_0_13_RW0_clk),
    .RW0_wdata(mem_0_13_RW0_wdata),
    .RW0_rdata(mem_0_13_RW0_rdata),
    .RW0_en(mem_0_13_RW0_en),
    .RW0_wmode(mem_0_13_RW0_wmode),
    .RW0_wmask(mem_0_13_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_14 (
    .RW0_addr(mem_0_14_RW0_addr),
    .RW0_clk(mem_0_14_RW0_clk),
    .RW0_wdata(mem_0_14_RW0_wdata),
    .RW0_rdata(mem_0_14_RW0_rdata),
    .RW0_en(mem_0_14_RW0_en),
    .RW0_wmode(mem_0_14_RW0_wmode),
    .RW0_wmask(mem_0_14_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_15 (
    .RW0_addr(mem_0_15_RW0_addr),
    .RW0_clk(mem_0_15_RW0_clk),
    .RW0_wdata(mem_0_15_RW0_wdata),
    .RW0_rdata(mem_0_15_RW0_rdata),
    .RW0_en(mem_0_15_RW0_en),
    .RW0_wmode(mem_0_15_RW0_wmode),
    .RW0_wmask(mem_0_15_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_16 (
    .RW0_addr(mem_0_16_RW0_addr),
    .RW0_clk(mem_0_16_RW0_clk),
    .RW0_wdata(mem_0_16_RW0_wdata),
    .RW0_rdata(mem_0_16_RW0_rdata),
    .RW0_en(mem_0_16_RW0_en),
    .RW0_wmode(mem_0_16_RW0_wmode),
    .RW0_wmask(mem_0_16_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_17 (
    .RW0_addr(mem_0_17_RW0_addr),
    .RW0_clk(mem_0_17_RW0_clk),
    .RW0_wdata(mem_0_17_RW0_wdata),
    .RW0_rdata(mem_0_17_RW0_rdata),
    .RW0_en(mem_0_17_RW0_en),
    .RW0_wmode(mem_0_17_RW0_wmode),
    .RW0_wmask(mem_0_17_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_18 (
    .RW0_addr(mem_0_18_RW0_addr),
    .RW0_clk(mem_0_18_RW0_clk),
    .RW0_wdata(mem_0_18_RW0_wdata),
    .RW0_rdata(mem_0_18_RW0_rdata),
    .RW0_en(mem_0_18_RW0_en),
    .RW0_wmode(mem_0_18_RW0_wmode),
    .RW0_wmask(mem_0_18_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_19 (
    .RW0_addr(mem_0_19_RW0_addr),
    .RW0_clk(mem_0_19_RW0_clk),
    .RW0_wdata(mem_0_19_RW0_wdata),
    .RW0_rdata(mem_0_19_RW0_rdata),
    .RW0_en(mem_0_19_RW0_en),
    .RW0_wmode(mem_0_19_RW0_wmode),
    .RW0_wmask(mem_0_19_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_20 (
    .RW0_addr(mem_0_20_RW0_addr),
    .RW0_clk(mem_0_20_RW0_clk),
    .RW0_wdata(mem_0_20_RW0_wdata),
    .RW0_rdata(mem_0_20_RW0_rdata),
    .RW0_en(mem_0_20_RW0_en),
    .RW0_wmode(mem_0_20_RW0_wmode),
    .RW0_wmask(mem_0_20_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_21 (
    .RW0_addr(mem_0_21_RW0_addr),
    .RW0_clk(mem_0_21_RW0_clk),
    .RW0_wdata(mem_0_21_RW0_wdata),
    .RW0_rdata(mem_0_21_RW0_rdata),
    .RW0_en(mem_0_21_RW0_en),
    .RW0_wmode(mem_0_21_RW0_wmode),
    .RW0_wmask(mem_0_21_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_22 (
    .RW0_addr(mem_0_22_RW0_addr),
    .RW0_clk(mem_0_22_RW0_clk),
    .RW0_wdata(mem_0_22_RW0_wdata),
    .RW0_rdata(mem_0_22_RW0_rdata),
    .RW0_en(mem_0_22_RW0_en),
    .RW0_wmode(mem_0_22_RW0_wmode),
    .RW0_wmask(mem_0_22_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_23 (
    .RW0_addr(mem_0_23_RW0_addr),
    .RW0_clk(mem_0_23_RW0_clk),
    .RW0_wdata(mem_0_23_RW0_wdata),
    .RW0_rdata(mem_0_23_RW0_rdata),
    .RW0_en(mem_0_23_RW0_en),
    .RW0_wmode(mem_0_23_RW0_wmode),
    .RW0_wmask(mem_0_23_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_24 (
    .RW0_addr(mem_0_24_RW0_addr),
    .RW0_clk(mem_0_24_RW0_clk),
    .RW0_wdata(mem_0_24_RW0_wdata),
    .RW0_rdata(mem_0_24_RW0_rdata),
    .RW0_en(mem_0_24_RW0_en),
    .RW0_wmode(mem_0_24_RW0_wmode),
    .RW0_wmask(mem_0_24_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_25 (
    .RW0_addr(mem_0_25_RW0_addr),
    .RW0_clk(mem_0_25_RW0_clk),
    .RW0_wdata(mem_0_25_RW0_wdata),
    .RW0_rdata(mem_0_25_RW0_rdata),
    .RW0_en(mem_0_25_RW0_en),
    .RW0_wmode(mem_0_25_RW0_wmode),
    .RW0_wmask(mem_0_25_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_26 (
    .RW0_addr(mem_0_26_RW0_addr),
    .RW0_clk(mem_0_26_RW0_clk),
    .RW0_wdata(mem_0_26_RW0_wdata),
    .RW0_rdata(mem_0_26_RW0_rdata),
    .RW0_en(mem_0_26_RW0_en),
    .RW0_wmode(mem_0_26_RW0_wmode),
    .RW0_wmask(mem_0_26_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_27 (
    .RW0_addr(mem_0_27_RW0_addr),
    .RW0_clk(mem_0_27_RW0_clk),
    .RW0_wdata(mem_0_27_RW0_wdata),
    .RW0_rdata(mem_0_27_RW0_rdata),
    .RW0_en(mem_0_27_RW0_en),
    .RW0_wmode(mem_0_27_RW0_wmode),
    .RW0_wmask(mem_0_27_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_28 (
    .RW0_addr(mem_0_28_RW0_addr),
    .RW0_clk(mem_0_28_RW0_clk),
    .RW0_wdata(mem_0_28_RW0_wdata),
    .RW0_rdata(mem_0_28_RW0_rdata),
    .RW0_en(mem_0_28_RW0_en),
    .RW0_wmode(mem_0_28_RW0_wmode),
    .RW0_wmask(mem_0_28_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_29 (
    .RW0_addr(mem_0_29_RW0_addr),
    .RW0_clk(mem_0_29_RW0_clk),
    .RW0_wdata(mem_0_29_RW0_wdata),
    .RW0_rdata(mem_0_29_RW0_rdata),
    .RW0_en(mem_0_29_RW0_en),
    .RW0_wmode(mem_0_29_RW0_wmode),
    .RW0_wmask(mem_0_29_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_30 (
    .RW0_addr(mem_0_30_RW0_addr),
    .RW0_clk(mem_0_30_RW0_clk),
    .RW0_wdata(mem_0_30_RW0_wdata),
    .RW0_rdata(mem_0_30_RW0_rdata),
    .RW0_en(mem_0_30_RW0_en),
    .RW0_wmode(mem_0_30_RW0_wmode),
    .RW0_wmask(mem_0_30_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_31 (
    .RW0_addr(mem_0_31_RW0_addr),
    .RW0_clk(mem_0_31_RW0_clk),
    .RW0_wdata(mem_0_31_RW0_wdata),
    .RW0_rdata(mem_0_31_RW0_rdata),
    .RW0_en(mem_0_31_RW0_en),
    .RW0_wmode(mem_0_31_RW0_wmode),
    .RW0_wmask(mem_0_31_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_31,_GEN_29};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_RW0_addr = RW0_addr;
  assign mem_0_4_RW0_clk = RW0_clk;
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32];
  assign mem_0_4_RW0_en = RW0_en;
  assign mem_0_4_RW0_wmode = RW0_wmode;
  assign mem_0_4_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_RW0_addr = RW0_addr;
  assign mem_0_5_RW0_clk = RW0_clk;
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40];
  assign mem_0_5_RW0_en = RW0_en;
  assign mem_0_5_RW0_wmode = RW0_wmode;
  assign mem_0_5_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_RW0_addr = RW0_addr;
  assign mem_0_6_RW0_clk = RW0_clk;
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48];
  assign mem_0_6_RW0_en = RW0_en;
  assign mem_0_6_RW0_wmode = RW0_wmode;
  assign mem_0_6_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_RW0_addr = RW0_addr;
  assign mem_0_7_RW0_clk = RW0_clk;
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56];
  assign mem_0_7_RW0_en = RW0_en;
  assign mem_0_7_RW0_wmode = RW0_wmode;
  assign mem_0_7_RW0_wmask = RW0_wmask[7];
  assign mem_0_8_RW0_addr = RW0_addr;
  assign mem_0_8_RW0_clk = RW0_clk;
  assign mem_0_8_RW0_wdata = RW0_wdata[71:64];
  assign mem_0_8_RW0_en = RW0_en;
  assign mem_0_8_RW0_wmode = RW0_wmode;
  assign mem_0_8_RW0_wmask = RW0_wmask[8];
  assign mem_0_9_RW0_addr = RW0_addr;
  assign mem_0_9_RW0_clk = RW0_clk;
  assign mem_0_9_RW0_wdata = RW0_wdata[79:72];
  assign mem_0_9_RW0_en = RW0_en;
  assign mem_0_9_RW0_wmode = RW0_wmode;
  assign mem_0_9_RW0_wmask = RW0_wmask[9];
  assign mem_0_10_RW0_addr = RW0_addr;
  assign mem_0_10_RW0_clk = RW0_clk;
  assign mem_0_10_RW0_wdata = RW0_wdata[87:80];
  assign mem_0_10_RW0_en = RW0_en;
  assign mem_0_10_RW0_wmode = RW0_wmode;
  assign mem_0_10_RW0_wmask = RW0_wmask[10];
  assign mem_0_11_RW0_addr = RW0_addr;
  assign mem_0_11_RW0_clk = RW0_clk;
  assign mem_0_11_RW0_wdata = RW0_wdata[95:88];
  assign mem_0_11_RW0_en = RW0_en;
  assign mem_0_11_RW0_wmode = RW0_wmode;
  assign mem_0_11_RW0_wmask = RW0_wmask[11];
  assign mem_0_12_RW0_addr = RW0_addr;
  assign mem_0_12_RW0_clk = RW0_clk;
  assign mem_0_12_RW0_wdata = RW0_wdata[103:96];
  assign mem_0_12_RW0_en = RW0_en;
  assign mem_0_12_RW0_wmode = RW0_wmode;
  assign mem_0_12_RW0_wmask = RW0_wmask[12];
  assign mem_0_13_RW0_addr = RW0_addr;
  assign mem_0_13_RW0_clk = RW0_clk;
  assign mem_0_13_RW0_wdata = RW0_wdata[111:104];
  assign mem_0_13_RW0_en = RW0_en;
  assign mem_0_13_RW0_wmode = RW0_wmode;
  assign mem_0_13_RW0_wmask = RW0_wmask[13];
  assign mem_0_14_RW0_addr = RW0_addr;
  assign mem_0_14_RW0_clk = RW0_clk;
  assign mem_0_14_RW0_wdata = RW0_wdata[119:112];
  assign mem_0_14_RW0_en = RW0_en;
  assign mem_0_14_RW0_wmode = RW0_wmode;
  assign mem_0_14_RW0_wmask = RW0_wmask[14];
  assign mem_0_15_RW0_addr = RW0_addr;
  assign mem_0_15_RW0_clk = RW0_clk;
  assign mem_0_15_RW0_wdata = RW0_wdata[127:120];
  assign mem_0_15_RW0_en = RW0_en;
  assign mem_0_15_RW0_wmode = RW0_wmode;
  assign mem_0_15_RW0_wmask = RW0_wmask[15];
  assign mem_0_16_RW0_addr = RW0_addr;
  assign mem_0_16_RW0_clk = RW0_clk;
  assign mem_0_16_RW0_wdata = RW0_wdata[135:128];
  assign mem_0_16_RW0_en = RW0_en;
  assign mem_0_16_RW0_wmode = RW0_wmode;
  assign mem_0_16_RW0_wmask = RW0_wmask[16];
  assign mem_0_17_RW0_addr = RW0_addr;
  assign mem_0_17_RW0_clk = RW0_clk;
  assign mem_0_17_RW0_wdata = RW0_wdata[143:136];
  assign mem_0_17_RW0_en = RW0_en;
  assign mem_0_17_RW0_wmode = RW0_wmode;
  assign mem_0_17_RW0_wmask = RW0_wmask[17];
  assign mem_0_18_RW0_addr = RW0_addr;
  assign mem_0_18_RW0_clk = RW0_clk;
  assign mem_0_18_RW0_wdata = RW0_wdata[151:144];
  assign mem_0_18_RW0_en = RW0_en;
  assign mem_0_18_RW0_wmode = RW0_wmode;
  assign mem_0_18_RW0_wmask = RW0_wmask[18];
  assign mem_0_19_RW0_addr = RW0_addr;
  assign mem_0_19_RW0_clk = RW0_clk;
  assign mem_0_19_RW0_wdata = RW0_wdata[159:152];
  assign mem_0_19_RW0_en = RW0_en;
  assign mem_0_19_RW0_wmode = RW0_wmode;
  assign mem_0_19_RW0_wmask = RW0_wmask[19];
  assign mem_0_20_RW0_addr = RW0_addr;
  assign mem_0_20_RW0_clk = RW0_clk;
  assign mem_0_20_RW0_wdata = RW0_wdata[167:160];
  assign mem_0_20_RW0_en = RW0_en;
  assign mem_0_20_RW0_wmode = RW0_wmode;
  assign mem_0_20_RW0_wmask = RW0_wmask[20];
  assign mem_0_21_RW0_addr = RW0_addr;
  assign mem_0_21_RW0_clk = RW0_clk;
  assign mem_0_21_RW0_wdata = RW0_wdata[175:168];
  assign mem_0_21_RW0_en = RW0_en;
  assign mem_0_21_RW0_wmode = RW0_wmode;
  assign mem_0_21_RW0_wmask = RW0_wmask[21];
  assign mem_0_22_RW0_addr = RW0_addr;
  assign mem_0_22_RW0_clk = RW0_clk;
  assign mem_0_22_RW0_wdata = RW0_wdata[183:176];
  assign mem_0_22_RW0_en = RW0_en;
  assign mem_0_22_RW0_wmode = RW0_wmode;
  assign mem_0_22_RW0_wmask = RW0_wmask[22];
  assign mem_0_23_RW0_addr = RW0_addr;
  assign mem_0_23_RW0_clk = RW0_clk;
  assign mem_0_23_RW0_wdata = RW0_wdata[191:184];
  assign mem_0_23_RW0_en = RW0_en;
  assign mem_0_23_RW0_wmode = RW0_wmode;
  assign mem_0_23_RW0_wmask = RW0_wmask[23];
  assign mem_0_24_RW0_addr = RW0_addr;
  assign mem_0_24_RW0_clk = RW0_clk;
  assign mem_0_24_RW0_wdata = RW0_wdata[199:192];
  assign mem_0_24_RW0_en = RW0_en;
  assign mem_0_24_RW0_wmode = RW0_wmode;
  assign mem_0_24_RW0_wmask = RW0_wmask[24];
  assign mem_0_25_RW0_addr = RW0_addr;
  assign mem_0_25_RW0_clk = RW0_clk;
  assign mem_0_25_RW0_wdata = RW0_wdata[207:200];
  assign mem_0_25_RW0_en = RW0_en;
  assign mem_0_25_RW0_wmode = RW0_wmode;
  assign mem_0_25_RW0_wmask = RW0_wmask[25];
  assign mem_0_26_RW0_addr = RW0_addr;
  assign mem_0_26_RW0_clk = RW0_clk;
  assign mem_0_26_RW0_wdata = RW0_wdata[215:208];
  assign mem_0_26_RW0_en = RW0_en;
  assign mem_0_26_RW0_wmode = RW0_wmode;
  assign mem_0_26_RW0_wmask = RW0_wmask[26];
  assign mem_0_27_RW0_addr = RW0_addr;
  assign mem_0_27_RW0_clk = RW0_clk;
  assign mem_0_27_RW0_wdata = RW0_wdata[223:216];
  assign mem_0_27_RW0_en = RW0_en;
  assign mem_0_27_RW0_wmode = RW0_wmode;
  assign mem_0_27_RW0_wmask = RW0_wmask[27];
  assign mem_0_28_RW0_addr = RW0_addr;
  assign mem_0_28_RW0_clk = RW0_clk;
  assign mem_0_28_RW0_wdata = RW0_wdata[231:224];
  assign mem_0_28_RW0_en = RW0_en;
  assign mem_0_28_RW0_wmode = RW0_wmode;
  assign mem_0_28_RW0_wmask = RW0_wmask[28];
  assign mem_0_29_RW0_addr = RW0_addr;
  assign mem_0_29_RW0_clk = RW0_clk;
  assign mem_0_29_RW0_wdata = RW0_wdata[239:232];
  assign mem_0_29_RW0_en = RW0_en;
  assign mem_0_29_RW0_wmode = RW0_wmode;
  assign mem_0_29_RW0_wmask = RW0_wmask[29];
  assign mem_0_30_RW0_addr = RW0_addr;
  assign mem_0_30_RW0_clk = RW0_clk;
  assign mem_0_30_RW0_wdata = RW0_wdata[247:240];
  assign mem_0_30_RW0_en = RW0_en;
  assign mem_0_30_RW0_wmode = RW0_wmode;
  assign mem_0_30_RW0_wmask = RW0_wmask[30];
  assign mem_0_31_RW0_addr = RW0_addr;
  assign mem_0_31_RW0_clk = RW0_clk;
  assign mem_0_31_RW0_wdata = RW0_wdata[255:248];
  assign mem_0_31_RW0_en = RW0_en;
  assign mem_0_31_RW0_wmode = RW0_wmode;
  assign mem_0_31_RW0_wmask = RW0_wmask[31];
endmodule
module tag_array_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [87:0] RW0_wdata,
  output [87:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [5:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [21:0] mem_0_0_RW0_wdata;
  wire [21:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [5:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [21:0] mem_0_1_RW0_wdata;
  wire [21:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [5:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [21:0] mem_0_2_RW0_wdata;
  wire [21:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [5:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [21:0] mem_0_3_RW0_wdata;
  wire [21:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [21:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [21:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [21:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [21:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [43:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [65:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [43:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [65:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_tag_array_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module mem_ext(
  input  [9:0]   W0_addr,
  input          W0_clk,
  input  [511:0] W0_data,
  input          W0_en,
  input  [63:0]  W0_mask,
  input  [9:0]   R0_addr,
  input          R0_clk,
  output [511:0] R0_data,
  input          R0_en
);
  wire [9:0] mem_0_0_W0_addr;
  wire  mem_0_0_W0_clk;
  wire [7:0] mem_0_0_W0_data;
  wire  mem_0_0_W0_en;
  wire  mem_0_0_W0_mask;
  wire [9:0] mem_0_0_R0_addr;
  wire  mem_0_0_R0_clk;
  wire [7:0] mem_0_0_R0_data;
  wire  mem_0_0_R0_en;
  wire [9:0] mem_0_1_W0_addr;
  wire  mem_0_1_W0_clk;
  wire [7:0] mem_0_1_W0_data;
  wire  mem_0_1_W0_en;
  wire  mem_0_1_W0_mask;
  wire [9:0] mem_0_1_R0_addr;
  wire  mem_0_1_R0_clk;
  wire [7:0] mem_0_1_R0_data;
  wire  mem_0_1_R0_en;
  wire [9:0] mem_0_2_W0_addr;
  wire  mem_0_2_W0_clk;
  wire [7:0] mem_0_2_W0_data;
  wire  mem_0_2_W0_en;
  wire  mem_0_2_W0_mask;
  wire [9:0] mem_0_2_R0_addr;
  wire  mem_0_2_R0_clk;
  wire [7:0] mem_0_2_R0_data;
  wire  mem_0_2_R0_en;
  wire [9:0] mem_0_3_W0_addr;
  wire  mem_0_3_W0_clk;
  wire [7:0] mem_0_3_W0_data;
  wire  mem_0_3_W0_en;
  wire  mem_0_3_W0_mask;
  wire [9:0] mem_0_3_R0_addr;
  wire  mem_0_3_R0_clk;
  wire [7:0] mem_0_3_R0_data;
  wire  mem_0_3_R0_en;
  wire [9:0] mem_0_4_W0_addr;
  wire  mem_0_4_W0_clk;
  wire [7:0] mem_0_4_W0_data;
  wire  mem_0_4_W0_en;
  wire  mem_0_4_W0_mask;
  wire [9:0] mem_0_4_R0_addr;
  wire  mem_0_4_R0_clk;
  wire [7:0] mem_0_4_R0_data;
  wire  mem_0_4_R0_en;
  wire [9:0] mem_0_5_W0_addr;
  wire  mem_0_5_W0_clk;
  wire [7:0] mem_0_5_W0_data;
  wire  mem_0_5_W0_en;
  wire  mem_0_5_W0_mask;
  wire [9:0] mem_0_5_R0_addr;
  wire  mem_0_5_R0_clk;
  wire [7:0] mem_0_5_R0_data;
  wire  mem_0_5_R0_en;
  wire [9:0] mem_0_6_W0_addr;
  wire  mem_0_6_W0_clk;
  wire [7:0] mem_0_6_W0_data;
  wire  mem_0_6_W0_en;
  wire  mem_0_6_W0_mask;
  wire [9:0] mem_0_6_R0_addr;
  wire  mem_0_6_R0_clk;
  wire [7:0] mem_0_6_R0_data;
  wire  mem_0_6_R0_en;
  wire [9:0] mem_0_7_W0_addr;
  wire  mem_0_7_W0_clk;
  wire [7:0] mem_0_7_W0_data;
  wire  mem_0_7_W0_en;
  wire  mem_0_7_W0_mask;
  wire [9:0] mem_0_7_R0_addr;
  wire  mem_0_7_R0_clk;
  wire [7:0] mem_0_7_R0_data;
  wire  mem_0_7_R0_en;
  wire [9:0] mem_0_8_W0_addr;
  wire  mem_0_8_W0_clk;
  wire [7:0] mem_0_8_W0_data;
  wire  mem_0_8_W0_en;
  wire  mem_0_8_W0_mask;
  wire [9:0] mem_0_8_R0_addr;
  wire  mem_0_8_R0_clk;
  wire [7:0] mem_0_8_R0_data;
  wire  mem_0_8_R0_en;
  wire [9:0] mem_0_9_W0_addr;
  wire  mem_0_9_W0_clk;
  wire [7:0] mem_0_9_W0_data;
  wire  mem_0_9_W0_en;
  wire  mem_0_9_W0_mask;
  wire [9:0] mem_0_9_R0_addr;
  wire  mem_0_9_R0_clk;
  wire [7:0] mem_0_9_R0_data;
  wire  mem_0_9_R0_en;
  wire [9:0] mem_0_10_W0_addr;
  wire  mem_0_10_W0_clk;
  wire [7:0] mem_0_10_W0_data;
  wire  mem_0_10_W0_en;
  wire  mem_0_10_W0_mask;
  wire [9:0] mem_0_10_R0_addr;
  wire  mem_0_10_R0_clk;
  wire [7:0] mem_0_10_R0_data;
  wire  mem_0_10_R0_en;
  wire [9:0] mem_0_11_W0_addr;
  wire  mem_0_11_W0_clk;
  wire [7:0] mem_0_11_W0_data;
  wire  mem_0_11_W0_en;
  wire  mem_0_11_W0_mask;
  wire [9:0] mem_0_11_R0_addr;
  wire  mem_0_11_R0_clk;
  wire [7:0] mem_0_11_R0_data;
  wire  mem_0_11_R0_en;
  wire [9:0] mem_0_12_W0_addr;
  wire  mem_0_12_W0_clk;
  wire [7:0] mem_0_12_W0_data;
  wire  mem_0_12_W0_en;
  wire  mem_0_12_W0_mask;
  wire [9:0] mem_0_12_R0_addr;
  wire  mem_0_12_R0_clk;
  wire [7:0] mem_0_12_R0_data;
  wire  mem_0_12_R0_en;
  wire [9:0] mem_0_13_W0_addr;
  wire  mem_0_13_W0_clk;
  wire [7:0] mem_0_13_W0_data;
  wire  mem_0_13_W0_en;
  wire  mem_0_13_W0_mask;
  wire [9:0] mem_0_13_R0_addr;
  wire  mem_0_13_R0_clk;
  wire [7:0] mem_0_13_R0_data;
  wire  mem_0_13_R0_en;
  wire [9:0] mem_0_14_W0_addr;
  wire  mem_0_14_W0_clk;
  wire [7:0] mem_0_14_W0_data;
  wire  mem_0_14_W0_en;
  wire  mem_0_14_W0_mask;
  wire [9:0] mem_0_14_R0_addr;
  wire  mem_0_14_R0_clk;
  wire [7:0] mem_0_14_R0_data;
  wire  mem_0_14_R0_en;
  wire [9:0] mem_0_15_W0_addr;
  wire  mem_0_15_W0_clk;
  wire [7:0] mem_0_15_W0_data;
  wire  mem_0_15_W0_en;
  wire  mem_0_15_W0_mask;
  wire [9:0] mem_0_15_R0_addr;
  wire  mem_0_15_R0_clk;
  wire [7:0] mem_0_15_R0_data;
  wire  mem_0_15_R0_en;
  wire [9:0] mem_0_16_W0_addr;
  wire  mem_0_16_W0_clk;
  wire [7:0] mem_0_16_W0_data;
  wire  mem_0_16_W0_en;
  wire  mem_0_16_W0_mask;
  wire [9:0] mem_0_16_R0_addr;
  wire  mem_0_16_R0_clk;
  wire [7:0] mem_0_16_R0_data;
  wire  mem_0_16_R0_en;
  wire [9:0] mem_0_17_W0_addr;
  wire  mem_0_17_W0_clk;
  wire [7:0] mem_0_17_W0_data;
  wire  mem_0_17_W0_en;
  wire  mem_0_17_W0_mask;
  wire [9:0] mem_0_17_R0_addr;
  wire  mem_0_17_R0_clk;
  wire [7:0] mem_0_17_R0_data;
  wire  mem_0_17_R0_en;
  wire [9:0] mem_0_18_W0_addr;
  wire  mem_0_18_W0_clk;
  wire [7:0] mem_0_18_W0_data;
  wire  mem_0_18_W0_en;
  wire  mem_0_18_W0_mask;
  wire [9:0] mem_0_18_R0_addr;
  wire  mem_0_18_R0_clk;
  wire [7:0] mem_0_18_R0_data;
  wire  mem_0_18_R0_en;
  wire [9:0] mem_0_19_W0_addr;
  wire  mem_0_19_W0_clk;
  wire [7:0] mem_0_19_W0_data;
  wire  mem_0_19_W0_en;
  wire  mem_0_19_W0_mask;
  wire [9:0] mem_0_19_R0_addr;
  wire  mem_0_19_R0_clk;
  wire [7:0] mem_0_19_R0_data;
  wire  mem_0_19_R0_en;
  wire [9:0] mem_0_20_W0_addr;
  wire  mem_0_20_W0_clk;
  wire [7:0] mem_0_20_W0_data;
  wire  mem_0_20_W0_en;
  wire  mem_0_20_W0_mask;
  wire [9:0] mem_0_20_R0_addr;
  wire  mem_0_20_R0_clk;
  wire [7:0] mem_0_20_R0_data;
  wire  mem_0_20_R0_en;
  wire [9:0] mem_0_21_W0_addr;
  wire  mem_0_21_W0_clk;
  wire [7:0] mem_0_21_W0_data;
  wire  mem_0_21_W0_en;
  wire  mem_0_21_W0_mask;
  wire [9:0] mem_0_21_R0_addr;
  wire  mem_0_21_R0_clk;
  wire [7:0] mem_0_21_R0_data;
  wire  mem_0_21_R0_en;
  wire [9:0] mem_0_22_W0_addr;
  wire  mem_0_22_W0_clk;
  wire [7:0] mem_0_22_W0_data;
  wire  mem_0_22_W0_en;
  wire  mem_0_22_W0_mask;
  wire [9:0] mem_0_22_R0_addr;
  wire  mem_0_22_R0_clk;
  wire [7:0] mem_0_22_R0_data;
  wire  mem_0_22_R0_en;
  wire [9:0] mem_0_23_W0_addr;
  wire  mem_0_23_W0_clk;
  wire [7:0] mem_0_23_W0_data;
  wire  mem_0_23_W0_en;
  wire  mem_0_23_W0_mask;
  wire [9:0] mem_0_23_R0_addr;
  wire  mem_0_23_R0_clk;
  wire [7:0] mem_0_23_R0_data;
  wire  mem_0_23_R0_en;
  wire [9:0] mem_0_24_W0_addr;
  wire  mem_0_24_W0_clk;
  wire [7:0] mem_0_24_W0_data;
  wire  mem_0_24_W0_en;
  wire  mem_0_24_W0_mask;
  wire [9:0] mem_0_24_R0_addr;
  wire  mem_0_24_R0_clk;
  wire [7:0] mem_0_24_R0_data;
  wire  mem_0_24_R0_en;
  wire [9:0] mem_0_25_W0_addr;
  wire  mem_0_25_W0_clk;
  wire [7:0] mem_0_25_W0_data;
  wire  mem_0_25_W0_en;
  wire  mem_0_25_W0_mask;
  wire [9:0] mem_0_25_R0_addr;
  wire  mem_0_25_R0_clk;
  wire [7:0] mem_0_25_R0_data;
  wire  mem_0_25_R0_en;
  wire [9:0] mem_0_26_W0_addr;
  wire  mem_0_26_W0_clk;
  wire [7:0] mem_0_26_W0_data;
  wire  mem_0_26_W0_en;
  wire  mem_0_26_W0_mask;
  wire [9:0] mem_0_26_R0_addr;
  wire  mem_0_26_R0_clk;
  wire [7:0] mem_0_26_R0_data;
  wire  mem_0_26_R0_en;
  wire [9:0] mem_0_27_W0_addr;
  wire  mem_0_27_W0_clk;
  wire [7:0] mem_0_27_W0_data;
  wire  mem_0_27_W0_en;
  wire  mem_0_27_W0_mask;
  wire [9:0] mem_0_27_R0_addr;
  wire  mem_0_27_R0_clk;
  wire [7:0] mem_0_27_R0_data;
  wire  mem_0_27_R0_en;
  wire [9:0] mem_0_28_W0_addr;
  wire  mem_0_28_W0_clk;
  wire [7:0] mem_0_28_W0_data;
  wire  mem_0_28_W0_en;
  wire  mem_0_28_W0_mask;
  wire [9:0] mem_0_28_R0_addr;
  wire  mem_0_28_R0_clk;
  wire [7:0] mem_0_28_R0_data;
  wire  mem_0_28_R0_en;
  wire [9:0] mem_0_29_W0_addr;
  wire  mem_0_29_W0_clk;
  wire [7:0] mem_0_29_W0_data;
  wire  mem_0_29_W0_en;
  wire  mem_0_29_W0_mask;
  wire [9:0] mem_0_29_R0_addr;
  wire  mem_0_29_R0_clk;
  wire [7:0] mem_0_29_R0_data;
  wire  mem_0_29_R0_en;
  wire [9:0] mem_0_30_W0_addr;
  wire  mem_0_30_W0_clk;
  wire [7:0] mem_0_30_W0_data;
  wire  mem_0_30_W0_en;
  wire  mem_0_30_W0_mask;
  wire [9:0] mem_0_30_R0_addr;
  wire  mem_0_30_R0_clk;
  wire [7:0] mem_0_30_R0_data;
  wire  mem_0_30_R0_en;
  wire [9:0] mem_0_31_W0_addr;
  wire  mem_0_31_W0_clk;
  wire [7:0] mem_0_31_W0_data;
  wire  mem_0_31_W0_en;
  wire  mem_0_31_W0_mask;
  wire [9:0] mem_0_31_R0_addr;
  wire  mem_0_31_R0_clk;
  wire [7:0] mem_0_31_R0_data;
  wire  mem_0_31_R0_en;
  wire [9:0] mem_0_32_W0_addr;
  wire  mem_0_32_W0_clk;
  wire [7:0] mem_0_32_W0_data;
  wire  mem_0_32_W0_en;
  wire  mem_0_32_W0_mask;
  wire [9:0] mem_0_32_R0_addr;
  wire  mem_0_32_R0_clk;
  wire [7:0] mem_0_32_R0_data;
  wire  mem_0_32_R0_en;
  wire [9:0] mem_0_33_W0_addr;
  wire  mem_0_33_W0_clk;
  wire [7:0] mem_0_33_W0_data;
  wire  mem_0_33_W0_en;
  wire  mem_0_33_W0_mask;
  wire [9:0] mem_0_33_R0_addr;
  wire  mem_0_33_R0_clk;
  wire [7:0] mem_0_33_R0_data;
  wire  mem_0_33_R0_en;
  wire [9:0] mem_0_34_W0_addr;
  wire  mem_0_34_W0_clk;
  wire [7:0] mem_0_34_W0_data;
  wire  mem_0_34_W0_en;
  wire  mem_0_34_W0_mask;
  wire [9:0] mem_0_34_R0_addr;
  wire  mem_0_34_R0_clk;
  wire [7:0] mem_0_34_R0_data;
  wire  mem_0_34_R0_en;
  wire [9:0] mem_0_35_W0_addr;
  wire  mem_0_35_W0_clk;
  wire [7:0] mem_0_35_W0_data;
  wire  mem_0_35_W0_en;
  wire  mem_0_35_W0_mask;
  wire [9:0] mem_0_35_R0_addr;
  wire  mem_0_35_R0_clk;
  wire [7:0] mem_0_35_R0_data;
  wire  mem_0_35_R0_en;
  wire [9:0] mem_0_36_W0_addr;
  wire  mem_0_36_W0_clk;
  wire [7:0] mem_0_36_W0_data;
  wire  mem_0_36_W0_en;
  wire  mem_0_36_W0_mask;
  wire [9:0] mem_0_36_R0_addr;
  wire  mem_0_36_R0_clk;
  wire [7:0] mem_0_36_R0_data;
  wire  mem_0_36_R0_en;
  wire [9:0] mem_0_37_W0_addr;
  wire  mem_0_37_W0_clk;
  wire [7:0] mem_0_37_W0_data;
  wire  mem_0_37_W0_en;
  wire  mem_0_37_W0_mask;
  wire [9:0] mem_0_37_R0_addr;
  wire  mem_0_37_R0_clk;
  wire [7:0] mem_0_37_R0_data;
  wire  mem_0_37_R0_en;
  wire [9:0] mem_0_38_W0_addr;
  wire  mem_0_38_W0_clk;
  wire [7:0] mem_0_38_W0_data;
  wire  mem_0_38_W0_en;
  wire  mem_0_38_W0_mask;
  wire [9:0] mem_0_38_R0_addr;
  wire  mem_0_38_R0_clk;
  wire [7:0] mem_0_38_R0_data;
  wire  mem_0_38_R0_en;
  wire [9:0] mem_0_39_W0_addr;
  wire  mem_0_39_W0_clk;
  wire [7:0] mem_0_39_W0_data;
  wire  mem_0_39_W0_en;
  wire  mem_0_39_W0_mask;
  wire [9:0] mem_0_39_R0_addr;
  wire  mem_0_39_R0_clk;
  wire [7:0] mem_0_39_R0_data;
  wire  mem_0_39_R0_en;
  wire [9:0] mem_0_40_W0_addr;
  wire  mem_0_40_W0_clk;
  wire [7:0] mem_0_40_W0_data;
  wire  mem_0_40_W0_en;
  wire  mem_0_40_W0_mask;
  wire [9:0] mem_0_40_R0_addr;
  wire  mem_0_40_R0_clk;
  wire [7:0] mem_0_40_R0_data;
  wire  mem_0_40_R0_en;
  wire [9:0] mem_0_41_W0_addr;
  wire  mem_0_41_W0_clk;
  wire [7:0] mem_0_41_W0_data;
  wire  mem_0_41_W0_en;
  wire  mem_0_41_W0_mask;
  wire [9:0] mem_0_41_R0_addr;
  wire  mem_0_41_R0_clk;
  wire [7:0] mem_0_41_R0_data;
  wire  mem_0_41_R0_en;
  wire [9:0] mem_0_42_W0_addr;
  wire  mem_0_42_W0_clk;
  wire [7:0] mem_0_42_W0_data;
  wire  mem_0_42_W0_en;
  wire  mem_0_42_W0_mask;
  wire [9:0] mem_0_42_R0_addr;
  wire  mem_0_42_R0_clk;
  wire [7:0] mem_0_42_R0_data;
  wire  mem_0_42_R0_en;
  wire [9:0] mem_0_43_W0_addr;
  wire  mem_0_43_W0_clk;
  wire [7:0] mem_0_43_W0_data;
  wire  mem_0_43_W0_en;
  wire  mem_0_43_W0_mask;
  wire [9:0] mem_0_43_R0_addr;
  wire  mem_0_43_R0_clk;
  wire [7:0] mem_0_43_R0_data;
  wire  mem_0_43_R0_en;
  wire [9:0] mem_0_44_W0_addr;
  wire  mem_0_44_W0_clk;
  wire [7:0] mem_0_44_W0_data;
  wire  mem_0_44_W0_en;
  wire  mem_0_44_W0_mask;
  wire [9:0] mem_0_44_R0_addr;
  wire  mem_0_44_R0_clk;
  wire [7:0] mem_0_44_R0_data;
  wire  mem_0_44_R0_en;
  wire [9:0] mem_0_45_W0_addr;
  wire  mem_0_45_W0_clk;
  wire [7:0] mem_0_45_W0_data;
  wire  mem_0_45_W0_en;
  wire  mem_0_45_W0_mask;
  wire [9:0] mem_0_45_R0_addr;
  wire  mem_0_45_R0_clk;
  wire [7:0] mem_0_45_R0_data;
  wire  mem_0_45_R0_en;
  wire [9:0] mem_0_46_W0_addr;
  wire  mem_0_46_W0_clk;
  wire [7:0] mem_0_46_W0_data;
  wire  mem_0_46_W0_en;
  wire  mem_0_46_W0_mask;
  wire [9:0] mem_0_46_R0_addr;
  wire  mem_0_46_R0_clk;
  wire [7:0] mem_0_46_R0_data;
  wire  mem_0_46_R0_en;
  wire [9:0] mem_0_47_W0_addr;
  wire  mem_0_47_W0_clk;
  wire [7:0] mem_0_47_W0_data;
  wire  mem_0_47_W0_en;
  wire  mem_0_47_W0_mask;
  wire [9:0] mem_0_47_R0_addr;
  wire  mem_0_47_R0_clk;
  wire [7:0] mem_0_47_R0_data;
  wire  mem_0_47_R0_en;
  wire [9:0] mem_0_48_W0_addr;
  wire  mem_0_48_W0_clk;
  wire [7:0] mem_0_48_W0_data;
  wire  mem_0_48_W0_en;
  wire  mem_0_48_W0_mask;
  wire [9:0] mem_0_48_R0_addr;
  wire  mem_0_48_R0_clk;
  wire [7:0] mem_0_48_R0_data;
  wire  mem_0_48_R0_en;
  wire [9:0] mem_0_49_W0_addr;
  wire  mem_0_49_W0_clk;
  wire [7:0] mem_0_49_W0_data;
  wire  mem_0_49_W0_en;
  wire  mem_0_49_W0_mask;
  wire [9:0] mem_0_49_R0_addr;
  wire  mem_0_49_R0_clk;
  wire [7:0] mem_0_49_R0_data;
  wire  mem_0_49_R0_en;
  wire [9:0] mem_0_50_W0_addr;
  wire  mem_0_50_W0_clk;
  wire [7:0] mem_0_50_W0_data;
  wire  mem_0_50_W0_en;
  wire  mem_0_50_W0_mask;
  wire [9:0] mem_0_50_R0_addr;
  wire  mem_0_50_R0_clk;
  wire [7:0] mem_0_50_R0_data;
  wire  mem_0_50_R0_en;
  wire [9:0] mem_0_51_W0_addr;
  wire  mem_0_51_W0_clk;
  wire [7:0] mem_0_51_W0_data;
  wire  mem_0_51_W0_en;
  wire  mem_0_51_W0_mask;
  wire [9:0] mem_0_51_R0_addr;
  wire  mem_0_51_R0_clk;
  wire [7:0] mem_0_51_R0_data;
  wire  mem_0_51_R0_en;
  wire [9:0] mem_0_52_W0_addr;
  wire  mem_0_52_W0_clk;
  wire [7:0] mem_0_52_W0_data;
  wire  mem_0_52_W0_en;
  wire  mem_0_52_W0_mask;
  wire [9:0] mem_0_52_R0_addr;
  wire  mem_0_52_R0_clk;
  wire [7:0] mem_0_52_R0_data;
  wire  mem_0_52_R0_en;
  wire [9:0] mem_0_53_W0_addr;
  wire  mem_0_53_W0_clk;
  wire [7:0] mem_0_53_W0_data;
  wire  mem_0_53_W0_en;
  wire  mem_0_53_W0_mask;
  wire [9:0] mem_0_53_R0_addr;
  wire  mem_0_53_R0_clk;
  wire [7:0] mem_0_53_R0_data;
  wire  mem_0_53_R0_en;
  wire [9:0] mem_0_54_W0_addr;
  wire  mem_0_54_W0_clk;
  wire [7:0] mem_0_54_W0_data;
  wire  mem_0_54_W0_en;
  wire  mem_0_54_W0_mask;
  wire [9:0] mem_0_54_R0_addr;
  wire  mem_0_54_R0_clk;
  wire [7:0] mem_0_54_R0_data;
  wire  mem_0_54_R0_en;
  wire [9:0] mem_0_55_W0_addr;
  wire  mem_0_55_W0_clk;
  wire [7:0] mem_0_55_W0_data;
  wire  mem_0_55_W0_en;
  wire  mem_0_55_W0_mask;
  wire [9:0] mem_0_55_R0_addr;
  wire  mem_0_55_R0_clk;
  wire [7:0] mem_0_55_R0_data;
  wire  mem_0_55_R0_en;
  wire [9:0] mem_0_56_W0_addr;
  wire  mem_0_56_W0_clk;
  wire [7:0] mem_0_56_W0_data;
  wire  mem_0_56_W0_en;
  wire  mem_0_56_W0_mask;
  wire [9:0] mem_0_56_R0_addr;
  wire  mem_0_56_R0_clk;
  wire [7:0] mem_0_56_R0_data;
  wire  mem_0_56_R0_en;
  wire [9:0] mem_0_57_W0_addr;
  wire  mem_0_57_W0_clk;
  wire [7:0] mem_0_57_W0_data;
  wire  mem_0_57_W0_en;
  wire  mem_0_57_W0_mask;
  wire [9:0] mem_0_57_R0_addr;
  wire  mem_0_57_R0_clk;
  wire [7:0] mem_0_57_R0_data;
  wire  mem_0_57_R0_en;
  wire [9:0] mem_0_58_W0_addr;
  wire  mem_0_58_W0_clk;
  wire [7:0] mem_0_58_W0_data;
  wire  mem_0_58_W0_en;
  wire  mem_0_58_W0_mask;
  wire [9:0] mem_0_58_R0_addr;
  wire  mem_0_58_R0_clk;
  wire [7:0] mem_0_58_R0_data;
  wire  mem_0_58_R0_en;
  wire [9:0] mem_0_59_W0_addr;
  wire  mem_0_59_W0_clk;
  wire [7:0] mem_0_59_W0_data;
  wire  mem_0_59_W0_en;
  wire  mem_0_59_W0_mask;
  wire [9:0] mem_0_59_R0_addr;
  wire  mem_0_59_R0_clk;
  wire [7:0] mem_0_59_R0_data;
  wire  mem_0_59_R0_en;
  wire [9:0] mem_0_60_W0_addr;
  wire  mem_0_60_W0_clk;
  wire [7:0] mem_0_60_W0_data;
  wire  mem_0_60_W0_en;
  wire  mem_0_60_W0_mask;
  wire [9:0] mem_0_60_R0_addr;
  wire  mem_0_60_R0_clk;
  wire [7:0] mem_0_60_R0_data;
  wire  mem_0_60_R0_en;
  wire [9:0] mem_0_61_W0_addr;
  wire  mem_0_61_W0_clk;
  wire [7:0] mem_0_61_W0_data;
  wire  mem_0_61_W0_en;
  wire  mem_0_61_W0_mask;
  wire [9:0] mem_0_61_R0_addr;
  wire  mem_0_61_R0_clk;
  wire [7:0] mem_0_61_R0_data;
  wire  mem_0_61_R0_en;
  wire [9:0] mem_0_62_W0_addr;
  wire  mem_0_62_W0_clk;
  wire [7:0] mem_0_62_W0_data;
  wire  mem_0_62_W0_en;
  wire  mem_0_62_W0_mask;
  wire [9:0] mem_0_62_R0_addr;
  wire  mem_0_62_R0_clk;
  wire [7:0] mem_0_62_R0_data;
  wire  mem_0_62_R0_en;
  wire [9:0] mem_0_63_W0_addr;
  wire  mem_0_63_W0_clk;
  wire [7:0] mem_0_63_W0_data;
  wire  mem_0_63_W0_en;
  wire  mem_0_63_W0_mask;
  wire [9:0] mem_0_63_R0_addr;
  wire  mem_0_63_R0_clk;
  wire [7:0] mem_0_63_R0_data;
  wire  mem_0_63_R0_en;
  wire [7:0] R0_data_0_0 = mem_0_0_R0_data;
  wire [7:0] R0_data_0_1 = mem_0_1_R0_data;
  wire [7:0] R0_data_0_2 = mem_0_2_R0_data;
  wire [7:0] R0_data_0_3 = mem_0_3_R0_data;
  wire [7:0] R0_data_0_4 = mem_0_4_R0_data;
  wire [7:0] R0_data_0_5 = mem_0_5_R0_data;
  wire [7:0] R0_data_0_6 = mem_0_6_R0_data;
  wire [7:0] R0_data_0_7 = mem_0_7_R0_data;
  wire [7:0] R0_data_0_8 = mem_0_8_R0_data;
  wire [7:0] R0_data_0_9 = mem_0_9_R0_data;
  wire [7:0] R0_data_0_10 = mem_0_10_R0_data;
  wire [7:0] R0_data_0_11 = mem_0_11_R0_data;
  wire [7:0] R0_data_0_12 = mem_0_12_R0_data;
  wire [7:0] R0_data_0_13 = mem_0_13_R0_data;
  wire [7:0] R0_data_0_14 = mem_0_14_R0_data;
  wire [7:0] R0_data_0_15 = mem_0_15_R0_data;
  wire [7:0] R0_data_0_16 = mem_0_16_R0_data;
  wire [7:0] R0_data_0_17 = mem_0_17_R0_data;
  wire [7:0] R0_data_0_18 = mem_0_18_R0_data;
  wire [7:0] R0_data_0_19 = mem_0_19_R0_data;
  wire [7:0] R0_data_0_20 = mem_0_20_R0_data;
  wire [7:0] R0_data_0_21 = mem_0_21_R0_data;
  wire [7:0] R0_data_0_22 = mem_0_22_R0_data;
  wire [7:0] R0_data_0_23 = mem_0_23_R0_data;
  wire [7:0] R0_data_0_24 = mem_0_24_R0_data;
  wire [7:0] R0_data_0_25 = mem_0_25_R0_data;
  wire [7:0] R0_data_0_26 = mem_0_26_R0_data;
  wire [7:0] R0_data_0_27 = mem_0_27_R0_data;
  wire [7:0] R0_data_0_28 = mem_0_28_R0_data;
  wire [7:0] R0_data_0_29 = mem_0_29_R0_data;
  wire [7:0] R0_data_0_30 = mem_0_30_R0_data;
  wire [7:0] R0_data_0_31 = mem_0_31_R0_data;
  wire [7:0] R0_data_0_32 = mem_0_32_R0_data;
  wire [7:0] R0_data_0_33 = mem_0_33_R0_data;
  wire [7:0] R0_data_0_34 = mem_0_34_R0_data;
  wire [7:0] R0_data_0_35 = mem_0_35_R0_data;
  wire [7:0] R0_data_0_36 = mem_0_36_R0_data;
  wire [7:0] R0_data_0_37 = mem_0_37_R0_data;
  wire [7:0] R0_data_0_38 = mem_0_38_R0_data;
  wire [7:0] R0_data_0_39 = mem_0_39_R0_data;
  wire [7:0] R0_data_0_40 = mem_0_40_R0_data;
  wire [7:0] R0_data_0_41 = mem_0_41_R0_data;
  wire [7:0] R0_data_0_42 = mem_0_42_R0_data;
  wire [7:0] R0_data_0_43 = mem_0_43_R0_data;
  wire [7:0] R0_data_0_44 = mem_0_44_R0_data;
  wire [7:0] R0_data_0_45 = mem_0_45_R0_data;
  wire [7:0] R0_data_0_46 = mem_0_46_R0_data;
  wire [7:0] R0_data_0_47 = mem_0_47_R0_data;
  wire [7:0] R0_data_0_48 = mem_0_48_R0_data;
  wire [7:0] R0_data_0_49 = mem_0_49_R0_data;
  wire [7:0] R0_data_0_50 = mem_0_50_R0_data;
  wire [7:0] R0_data_0_51 = mem_0_51_R0_data;
  wire [7:0] R0_data_0_52 = mem_0_52_R0_data;
  wire [7:0] R0_data_0_53 = mem_0_53_R0_data;
  wire [7:0] R0_data_0_54 = mem_0_54_R0_data;
  wire [7:0] R0_data_0_55 = mem_0_55_R0_data;
  wire [7:0] R0_data_0_56 = mem_0_56_R0_data;
  wire [7:0] R0_data_0_57 = mem_0_57_R0_data;
  wire [7:0] R0_data_0_58 = mem_0_58_R0_data;
  wire [7:0] R0_data_0_59 = mem_0_59_R0_data;
  wire [7:0] R0_data_0_60 = mem_0_60_R0_data;
  wire [7:0] R0_data_0_61 = mem_0_61_R0_data;
  wire [7:0] R0_data_0_62 = mem_0_62_R0_data;
  wire [7:0] R0_data_0_63 = mem_0_63_R0_data;
  wire [15:0] _GEN_0 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_2 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_3 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_4 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_5 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_6 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}
    ;
  wire [71:0] _GEN_7 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,
    R0_data_0_0};
  wire [79:0] _GEN_8 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,
    R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_9 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_14 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_15 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_16 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_17 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_18 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_19 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_20 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_21 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_22 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_23 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_24 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_25 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_26 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_27 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_28 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_29 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_30 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_31 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_32 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_33 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_34 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_35 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_36 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_37 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_38 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_39 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_40 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_41 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_42 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_43 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_44 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_45 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_46 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_47 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_48 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_49 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_50 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_51 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_52 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_53 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_54 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_55 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_56 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_57 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_58 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_59 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_60 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_61 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  wire [511:0] R0_data_0 = {R0_data_0_63,R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,
    R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [15:0] _GEN_62 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_63 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_64 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_65 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_66 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_67 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_68 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0
    };
  wire [71:0] _GEN_69 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1
    ,R0_data_0_0};
  wire [79:0] _GEN_70 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2
    ,R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_71 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_72 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_73 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_74 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_75 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_76 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_77 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_78 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_79 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_80 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_81 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_82 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_83 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_84 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_85 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_86 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_87 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_88 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_89 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_90 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_91 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_92 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_93 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_94 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_95 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_96 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_97 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_98 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_99 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_100 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_101 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_102 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_103 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_104 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_105 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_106 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_107 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_108 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_109 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_110 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_111 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_112 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_113 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_114 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_115 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_116 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_117 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_118 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_119 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_120 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_121 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_122 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_123 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  split_mem_ext mem_0_0 (
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_mem_ext mem_0_1 (
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_mem_ext mem_0_2 (
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_mem_ext mem_0_3 (
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  split_mem_ext mem_0_4 (
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask),
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en)
  );
  split_mem_ext mem_0_5 (
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask),
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en)
  );
  split_mem_ext mem_0_6 (
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask),
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en)
  );
  split_mem_ext mem_0_7 (
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask),
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en)
  );
  split_mem_ext mem_0_8 (
    .W0_addr(mem_0_8_W0_addr),
    .W0_clk(mem_0_8_W0_clk),
    .W0_data(mem_0_8_W0_data),
    .W0_en(mem_0_8_W0_en),
    .W0_mask(mem_0_8_W0_mask),
    .R0_addr(mem_0_8_R0_addr),
    .R0_clk(mem_0_8_R0_clk),
    .R0_data(mem_0_8_R0_data),
    .R0_en(mem_0_8_R0_en)
  );
  split_mem_ext mem_0_9 (
    .W0_addr(mem_0_9_W0_addr),
    .W0_clk(mem_0_9_W0_clk),
    .W0_data(mem_0_9_W0_data),
    .W0_en(mem_0_9_W0_en),
    .W0_mask(mem_0_9_W0_mask),
    .R0_addr(mem_0_9_R0_addr),
    .R0_clk(mem_0_9_R0_clk),
    .R0_data(mem_0_9_R0_data),
    .R0_en(mem_0_9_R0_en)
  );
  split_mem_ext mem_0_10 (
    .W0_addr(mem_0_10_W0_addr),
    .W0_clk(mem_0_10_W0_clk),
    .W0_data(mem_0_10_W0_data),
    .W0_en(mem_0_10_W0_en),
    .W0_mask(mem_0_10_W0_mask),
    .R0_addr(mem_0_10_R0_addr),
    .R0_clk(mem_0_10_R0_clk),
    .R0_data(mem_0_10_R0_data),
    .R0_en(mem_0_10_R0_en)
  );
  split_mem_ext mem_0_11 (
    .W0_addr(mem_0_11_W0_addr),
    .W0_clk(mem_0_11_W0_clk),
    .W0_data(mem_0_11_W0_data),
    .W0_en(mem_0_11_W0_en),
    .W0_mask(mem_0_11_W0_mask),
    .R0_addr(mem_0_11_R0_addr),
    .R0_clk(mem_0_11_R0_clk),
    .R0_data(mem_0_11_R0_data),
    .R0_en(mem_0_11_R0_en)
  );
  split_mem_ext mem_0_12 (
    .W0_addr(mem_0_12_W0_addr),
    .W0_clk(mem_0_12_W0_clk),
    .W0_data(mem_0_12_W0_data),
    .W0_en(mem_0_12_W0_en),
    .W0_mask(mem_0_12_W0_mask),
    .R0_addr(mem_0_12_R0_addr),
    .R0_clk(mem_0_12_R0_clk),
    .R0_data(mem_0_12_R0_data),
    .R0_en(mem_0_12_R0_en)
  );
  split_mem_ext mem_0_13 (
    .W0_addr(mem_0_13_W0_addr),
    .W0_clk(mem_0_13_W0_clk),
    .W0_data(mem_0_13_W0_data),
    .W0_en(mem_0_13_W0_en),
    .W0_mask(mem_0_13_W0_mask),
    .R0_addr(mem_0_13_R0_addr),
    .R0_clk(mem_0_13_R0_clk),
    .R0_data(mem_0_13_R0_data),
    .R0_en(mem_0_13_R0_en)
  );
  split_mem_ext mem_0_14 (
    .W0_addr(mem_0_14_W0_addr),
    .W0_clk(mem_0_14_W0_clk),
    .W0_data(mem_0_14_W0_data),
    .W0_en(mem_0_14_W0_en),
    .W0_mask(mem_0_14_W0_mask),
    .R0_addr(mem_0_14_R0_addr),
    .R0_clk(mem_0_14_R0_clk),
    .R0_data(mem_0_14_R0_data),
    .R0_en(mem_0_14_R0_en)
  );
  split_mem_ext mem_0_15 (
    .W0_addr(mem_0_15_W0_addr),
    .W0_clk(mem_0_15_W0_clk),
    .W0_data(mem_0_15_W0_data),
    .W0_en(mem_0_15_W0_en),
    .W0_mask(mem_0_15_W0_mask),
    .R0_addr(mem_0_15_R0_addr),
    .R0_clk(mem_0_15_R0_clk),
    .R0_data(mem_0_15_R0_data),
    .R0_en(mem_0_15_R0_en)
  );
  split_mem_ext mem_0_16 (
    .W0_addr(mem_0_16_W0_addr),
    .W0_clk(mem_0_16_W0_clk),
    .W0_data(mem_0_16_W0_data),
    .W0_en(mem_0_16_W0_en),
    .W0_mask(mem_0_16_W0_mask),
    .R0_addr(mem_0_16_R0_addr),
    .R0_clk(mem_0_16_R0_clk),
    .R0_data(mem_0_16_R0_data),
    .R0_en(mem_0_16_R0_en)
  );
  split_mem_ext mem_0_17 (
    .W0_addr(mem_0_17_W0_addr),
    .W0_clk(mem_0_17_W0_clk),
    .W0_data(mem_0_17_W0_data),
    .W0_en(mem_0_17_W0_en),
    .W0_mask(mem_0_17_W0_mask),
    .R0_addr(mem_0_17_R0_addr),
    .R0_clk(mem_0_17_R0_clk),
    .R0_data(mem_0_17_R0_data),
    .R0_en(mem_0_17_R0_en)
  );
  split_mem_ext mem_0_18 (
    .W0_addr(mem_0_18_W0_addr),
    .W0_clk(mem_0_18_W0_clk),
    .W0_data(mem_0_18_W0_data),
    .W0_en(mem_0_18_W0_en),
    .W0_mask(mem_0_18_W0_mask),
    .R0_addr(mem_0_18_R0_addr),
    .R0_clk(mem_0_18_R0_clk),
    .R0_data(mem_0_18_R0_data),
    .R0_en(mem_0_18_R0_en)
  );
  split_mem_ext mem_0_19 (
    .W0_addr(mem_0_19_W0_addr),
    .W0_clk(mem_0_19_W0_clk),
    .W0_data(mem_0_19_W0_data),
    .W0_en(mem_0_19_W0_en),
    .W0_mask(mem_0_19_W0_mask),
    .R0_addr(mem_0_19_R0_addr),
    .R0_clk(mem_0_19_R0_clk),
    .R0_data(mem_0_19_R0_data),
    .R0_en(mem_0_19_R0_en)
  );
  split_mem_ext mem_0_20 (
    .W0_addr(mem_0_20_W0_addr),
    .W0_clk(mem_0_20_W0_clk),
    .W0_data(mem_0_20_W0_data),
    .W0_en(mem_0_20_W0_en),
    .W0_mask(mem_0_20_W0_mask),
    .R0_addr(mem_0_20_R0_addr),
    .R0_clk(mem_0_20_R0_clk),
    .R0_data(mem_0_20_R0_data),
    .R0_en(mem_0_20_R0_en)
  );
  split_mem_ext mem_0_21 (
    .W0_addr(mem_0_21_W0_addr),
    .W0_clk(mem_0_21_W0_clk),
    .W0_data(mem_0_21_W0_data),
    .W0_en(mem_0_21_W0_en),
    .W0_mask(mem_0_21_W0_mask),
    .R0_addr(mem_0_21_R0_addr),
    .R0_clk(mem_0_21_R0_clk),
    .R0_data(mem_0_21_R0_data),
    .R0_en(mem_0_21_R0_en)
  );
  split_mem_ext mem_0_22 (
    .W0_addr(mem_0_22_W0_addr),
    .W0_clk(mem_0_22_W0_clk),
    .W0_data(mem_0_22_W0_data),
    .W0_en(mem_0_22_W0_en),
    .W0_mask(mem_0_22_W0_mask),
    .R0_addr(mem_0_22_R0_addr),
    .R0_clk(mem_0_22_R0_clk),
    .R0_data(mem_0_22_R0_data),
    .R0_en(mem_0_22_R0_en)
  );
  split_mem_ext mem_0_23 (
    .W0_addr(mem_0_23_W0_addr),
    .W0_clk(mem_0_23_W0_clk),
    .W0_data(mem_0_23_W0_data),
    .W0_en(mem_0_23_W0_en),
    .W0_mask(mem_0_23_W0_mask),
    .R0_addr(mem_0_23_R0_addr),
    .R0_clk(mem_0_23_R0_clk),
    .R0_data(mem_0_23_R0_data),
    .R0_en(mem_0_23_R0_en)
  );
  split_mem_ext mem_0_24 (
    .W0_addr(mem_0_24_W0_addr),
    .W0_clk(mem_0_24_W0_clk),
    .W0_data(mem_0_24_W0_data),
    .W0_en(mem_0_24_W0_en),
    .W0_mask(mem_0_24_W0_mask),
    .R0_addr(mem_0_24_R0_addr),
    .R0_clk(mem_0_24_R0_clk),
    .R0_data(mem_0_24_R0_data),
    .R0_en(mem_0_24_R0_en)
  );
  split_mem_ext mem_0_25 (
    .W0_addr(mem_0_25_W0_addr),
    .W0_clk(mem_0_25_W0_clk),
    .W0_data(mem_0_25_W0_data),
    .W0_en(mem_0_25_W0_en),
    .W0_mask(mem_0_25_W0_mask),
    .R0_addr(mem_0_25_R0_addr),
    .R0_clk(mem_0_25_R0_clk),
    .R0_data(mem_0_25_R0_data),
    .R0_en(mem_0_25_R0_en)
  );
  split_mem_ext mem_0_26 (
    .W0_addr(mem_0_26_W0_addr),
    .W0_clk(mem_0_26_W0_clk),
    .W0_data(mem_0_26_W0_data),
    .W0_en(mem_0_26_W0_en),
    .W0_mask(mem_0_26_W0_mask),
    .R0_addr(mem_0_26_R0_addr),
    .R0_clk(mem_0_26_R0_clk),
    .R0_data(mem_0_26_R0_data),
    .R0_en(mem_0_26_R0_en)
  );
  split_mem_ext mem_0_27 (
    .W0_addr(mem_0_27_W0_addr),
    .W0_clk(mem_0_27_W0_clk),
    .W0_data(mem_0_27_W0_data),
    .W0_en(mem_0_27_W0_en),
    .W0_mask(mem_0_27_W0_mask),
    .R0_addr(mem_0_27_R0_addr),
    .R0_clk(mem_0_27_R0_clk),
    .R0_data(mem_0_27_R0_data),
    .R0_en(mem_0_27_R0_en)
  );
  split_mem_ext mem_0_28 (
    .W0_addr(mem_0_28_W0_addr),
    .W0_clk(mem_0_28_W0_clk),
    .W0_data(mem_0_28_W0_data),
    .W0_en(mem_0_28_W0_en),
    .W0_mask(mem_0_28_W0_mask),
    .R0_addr(mem_0_28_R0_addr),
    .R0_clk(mem_0_28_R0_clk),
    .R0_data(mem_0_28_R0_data),
    .R0_en(mem_0_28_R0_en)
  );
  split_mem_ext mem_0_29 (
    .W0_addr(mem_0_29_W0_addr),
    .W0_clk(mem_0_29_W0_clk),
    .W0_data(mem_0_29_W0_data),
    .W0_en(mem_0_29_W0_en),
    .W0_mask(mem_0_29_W0_mask),
    .R0_addr(mem_0_29_R0_addr),
    .R0_clk(mem_0_29_R0_clk),
    .R0_data(mem_0_29_R0_data),
    .R0_en(mem_0_29_R0_en)
  );
  split_mem_ext mem_0_30 (
    .W0_addr(mem_0_30_W0_addr),
    .W0_clk(mem_0_30_W0_clk),
    .W0_data(mem_0_30_W0_data),
    .W0_en(mem_0_30_W0_en),
    .W0_mask(mem_0_30_W0_mask),
    .R0_addr(mem_0_30_R0_addr),
    .R0_clk(mem_0_30_R0_clk),
    .R0_data(mem_0_30_R0_data),
    .R0_en(mem_0_30_R0_en)
  );
  split_mem_ext mem_0_31 (
    .W0_addr(mem_0_31_W0_addr),
    .W0_clk(mem_0_31_W0_clk),
    .W0_data(mem_0_31_W0_data),
    .W0_en(mem_0_31_W0_en),
    .W0_mask(mem_0_31_W0_mask),
    .R0_addr(mem_0_31_R0_addr),
    .R0_clk(mem_0_31_R0_clk),
    .R0_data(mem_0_31_R0_data),
    .R0_en(mem_0_31_R0_en)
  );
  split_mem_ext mem_0_32 (
    .W0_addr(mem_0_32_W0_addr),
    .W0_clk(mem_0_32_W0_clk),
    .W0_data(mem_0_32_W0_data),
    .W0_en(mem_0_32_W0_en),
    .W0_mask(mem_0_32_W0_mask),
    .R0_addr(mem_0_32_R0_addr),
    .R0_clk(mem_0_32_R0_clk),
    .R0_data(mem_0_32_R0_data),
    .R0_en(mem_0_32_R0_en)
  );
  split_mem_ext mem_0_33 (
    .W0_addr(mem_0_33_W0_addr),
    .W0_clk(mem_0_33_W0_clk),
    .W0_data(mem_0_33_W0_data),
    .W0_en(mem_0_33_W0_en),
    .W0_mask(mem_0_33_W0_mask),
    .R0_addr(mem_0_33_R0_addr),
    .R0_clk(mem_0_33_R0_clk),
    .R0_data(mem_0_33_R0_data),
    .R0_en(mem_0_33_R0_en)
  );
  split_mem_ext mem_0_34 (
    .W0_addr(mem_0_34_W0_addr),
    .W0_clk(mem_0_34_W0_clk),
    .W0_data(mem_0_34_W0_data),
    .W0_en(mem_0_34_W0_en),
    .W0_mask(mem_0_34_W0_mask),
    .R0_addr(mem_0_34_R0_addr),
    .R0_clk(mem_0_34_R0_clk),
    .R0_data(mem_0_34_R0_data),
    .R0_en(mem_0_34_R0_en)
  );
  split_mem_ext mem_0_35 (
    .W0_addr(mem_0_35_W0_addr),
    .W0_clk(mem_0_35_W0_clk),
    .W0_data(mem_0_35_W0_data),
    .W0_en(mem_0_35_W0_en),
    .W0_mask(mem_0_35_W0_mask),
    .R0_addr(mem_0_35_R0_addr),
    .R0_clk(mem_0_35_R0_clk),
    .R0_data(mem_0_35_R0_data),
    .R0_en(mem_0_35_R0_en)
  );
  split_mem_ext mem_0_36 (
    .W0_addr(mem_0_36_W0_addr),
    .W0_clk(mem_0_36_W0_clk),
    .W0_data(mem_0_36_W0_data),
    .W0_en(mem_0_36_W0_en),
    .W0_mask(mem_0_36_W0_mask),
    .R0_addr(mem_0_36_R0_addr),
    .R0_clk(mem_0_36_R0_clk),
    .R0_data(mem_0_36_R0_data),
    .R0_en(mem_0_36_R0_en)
  );
  split_mem_ext mem_0_37 (
    .W0_addr(mem_0_37_W0_addr),
    .W0_clk(mem_0_37_W0_clk),
    .W0_data(mem_0_37_W0_data),
    .W0_en(mem_0_37_W0_en),
    .W0_mask(mem_0_37_W0_mask),
    .R0_addr(mem_0_37_R0_addr),
    .R0_clk(mem_0_37_R0_clk),
    .R0_data(mem_0_37_R0_data),
    .R0_en(mem_0_37_R0_en)
  );
  split_mem_ext mem_0_38 (
    .W0_addr(mem_0_38_W0_addr),
    .W0_clk(mem_0_38_W0_clk),
    .W0_data(mem_0_38_W0_data),
    .W0_en(mem_0_38_W0_en),
    .W0_mask(mem_0_38_W0_mask),
    .R0_addr(mem_0_38_R0_addr),
    .R0_clk(mem_0_38_R0_clk),
    .R0_data(mem_0_38_R0_data),
    .R0_en(mem_0_38_R0_en)
  );
  split_mem_ext mem_0_39 (
    .W0_addr(mem_0_39_W0_addr),
    .W0_clk(mem_0_39_W0_clk),
    .W0_data(mem_0_39_W0_data),
    .W0_en(mem_0_39_W0_en),
    .W0_mask(mem_0_39_W0_mask),
    .R0_addr(mem_0_39_R0_addr),
    .R0_clk(mem_0_39_R0_clk),
    .R0_data(mem_0_39_R0_data),
    .R0_en(mem_0_39_R0_en)
  );
  split_mem_ext mem_0_40 (
    .W0_addr(mem_0_40_W0_addr),
    .W0_clk(mem_0_40_W0_clk),
    .W0_data(mem_0_40_W0_data),
    .W0_en(mem_0_40_W0_en),
    .W0_mask(mem_0_40_W0_mask),
    .R0_addr(mem_0_40_R0_addr),
    .R0_clk(mem_0_40_R0_clk),
    .R0_data(mem_0_40_R0_data),
    .R0_en(mem_0_40_R0_en)
  );
  split_mem_ext mem_0_41 (
    .W0_addr(mem_0_41_W0_addr),
    .W0_clk(mem_0_41_W0_clk),
    .W0_data(mem_0_41_W0_data),
    .W0_en(mem_0_41_W0_en),
    .W0_mask(mem_0_41_W0_mask),
    .R0_addr(mem_0_41_R0_addr),
    .R0_clk(mem_0_41_R0_clk),
    .R0_data(mem_0_41_R0_data),
    .R0_en(mem_0_41_R0_en)
  );
  split_mem_ext mem_0_42 (
    .W0_addr(mem_0_42_W0_addr),
    .W0_clk(mem_0_42_W0_clk),
    .W0_data(mem_0_42_W0_data),
    .W0_en(mem_0_42_W0_en),
    .W0_mask(mem_0_42_W0_mask),
    .R0_addr(mem_0_42_R0_addr),
    .R0_clk(mem_0_42_R0_clk),
    .R0_data(mem_0_42_R0_data),
    .R0_en(mem_0_42_R0_en)
  );
  split_mem_ext mem_0_43 (
    .W0_addr(mem_0_43_W0_addr),
    .W0_clk(mem_0_43_W0_clk),
    .W0_data(mem_0_43_W0_data),
    .W0_en(mem_0_43_W0_en),
    .W0_mask(mem_0_43_W0_mask),
    .R0_addr(mem_0_43_R0_addr),
    .R0_clk(mem_0_43_R0_clk),
    .R0_data(mem_0_43_R0_data),
    .R0_en(mem_0_43_R0_en)
  );
  split_mem_ext mem_0_44 (
    .W0_addr(mem_0_44_W0_addr),
    .W0_clk(mem_0_44_W0_clk),
    .W0_data(mem_0_44_W0_data),
    .W0_en(mem_0_44_W0_en),
    .W0_mask(mem_0_44_W0_mask),
    .R0_addr(mem_0_44_R0_addr),
    .R0_clk(mem_0_44_R0_clk),
    .R0_data(mem_0_44_R0_data),
    .R0_en(mem_0_44_R0_en)
  );
  split_mem_ext mem_0_45 (
    .W0_addr(mem_0_45_W0_addr),
    .W0_clk(mem_0_45_W0_clk),
    .W0_data(mem_0_45_W0_data),
    .W0_en(mem_0_45_W0_en),
    .W0_mask(mem_0_45_W0_mask),
    .R0_addr(mem_0_45_R0_addr),
    .R0_clk(mem_0_45_R0_clk),
    .R0_data(mem_0_45_R0_data),
    .R0_en(mem_0_45_R0_en)
  );
  split_mem_ext mem_0_46 (
    .W0_addr(mem_0_46_W0_addr),
    .W0_clk(mem_0_46_W0_clk),
    .W0_data(mem_0_46_W0_data),
    .W0_en(mem_0_46_W0_en),
    .W0_mask(mem_0_46_W0_mask),
    .R0_addr(mem_0_46_R0_addr),
    .R0_clk(mem_0_46_R0_clk),
    .R0_data(mem_0_46_R0_data),
    .R0_en(mem_0_46_R0_en)
  );
  split_mem_ext mem_0_47 (
    .W0_addr(mem_0_47_W0_addr),
    .W0_clk(mem_0_47_W0_clk),
    .W0_data(mem_0_47_W0_data),
    .W0_en(mem_0_47_W0_en),
    .W0_mask(mem_0_47_W0_mask),
    .R0_addr(mem_0_47_R0_addr),
    .R0_clk(mem_0_47_R0_clk),
    .R0_data(mem_0_47_R0_data),
    .R0_en(mem_0_47_R0_en)
  );
  split_mem_ext mem_0_48 (
    .W0_addr(mem_0_48_W0_addr),
    .W0_clk(mem_0_48_W0_clk),
    .W0_data(mem_0_48_W0_data),
    .W0_en(mem_0_48_W0_en),
    .W0_mask(mem_0_48_W0_mask),
    .R0_addr(mem_0_48_R0_addr),
    .R0_clk(mem_0_48_R0_clk),
    .R0_data(mem_0_48_R0_data),
    .R0_en(mem_0_48_R0_en)
  );
  split_mem_ext mem_0_49 (
    .W0_addr(mem_0_49_W0_addr),
    .W0_clk(mem_0_49_W0_clk),
    .W0_data(mem_0_49_W0_data),
    .W0_en(mem_0_49_W0_en),
    .W0_mask(mem_0_49_W0_mask),
    .R0_addr(mem_0_49_R0_addr),
    .R0_clk(mem_0_49_R0_clk),
    .R0_data(mem_0_49_R0_data),
    .R0_en(mem_0_49_R0_en)
  );
  split_mem_ext mem_0_50 (
    .W0_addr(mem_0_50_W0_addr),
    .W0_clk(mem_0_50_W0_clk),
    .W0_data(mem_0_50_W0_data),
    .W0_en(mem_0_50_W0_en),
    .W0_mask(mem_0_50_W0_mask),
    .R0_addr(mem_0_50_R0_addr),
    .R0_clk(mem_0_50_R0_clk),
    .R0_data(mem_0_50_R0_data),
    .R0_en(mem_0_50_R0_en)
  );
  split_mem_ext mem_0_51 (
    .W0_addr(mem_0_51_W0_addr),
    .W0_clk(mem_0_51_W0_clk),
    .W0_data(mem_0_51_W0_data),
    .W0_en(mem_0_51_W0_en),
    .W0_mask(mem_0_51_W0_mask),
    .R0_addr(mem_0_51_R0_addr),
    .R0_clk(mem_0_51_R0_clk),
    .R0_data(mem_0_51_R0_data),
    .R0_en(mem_0_51_R0_en)
  );
  split_mem_ext mem_0_52 (
    .W0_addr(mem_0_52_W0_addr),
    .W0_clk(mem_0_52_W0_clk),
    .W0_data(mem_0_52_W0_data),
    .W0_en(mem_0_52_W0_en),
    .W0_mask(mem_0_52_W0_mask),
    .R0_addr(mem_0_52_R0_addr),
    .R0_clk(mem_0_52_R0_clk),
    .R0_data(mem_0_52_R0_data),
    .R0_en(mem_0_52_R0_en)
  );
  split_mem_ext mem_0_53 (
    .W0_addr(mem_0_53_W0_addr),
    .W0_clk(mem_0_53_W0_clk),
    .W0_data(mem_0_53_W0_data),
    .W0_en(mem_0_53_W0_en),
    .W0_mask(mem_0_53_W0_mask),
    .R0_addr(mem_0_53_R0_addr),
    .R0_clk(mem_0_53_R0_clk),
    .R0_data(mem_0_53_R0_data),
    .R0_en(mem_0_53_R0_en)
  );
  split_mem_ext mem_0_54 (
    .W0_addr(mem_0_54_W0_addr),
    .W0_clk(mem_0_54_W0_clk),
    .W0_data(mem_0_54_W0_data),
    .W0_en(mem_0_54_W0_en),
    .W0_mask(mem_0_54_W0_mask),
    .R0_addr(mem_0_54_R0_addr),
    .R0_clk(mem_0_54_R0_clk),
    .R0_data(mem_0_54_R0_data),
    .R0_en(mem_0_54_R0_en)
  );
  split_mem_ext mem_0_55 (
    .W0_addr(mem_0_55_W0_addr),
    .W0_clk(mem_0_55_W0_clk),
    .W0_data(mem_0_55_W0_data),
    .W0_en(mem_0_55_W0_en),
    .W0_mask(mem_0_55_W0_mask),
    .R0_addr(mem_0_55_R0_addr),
    .R0_clk(mem_0_55_R0_clk),
    .R0_data(mem_0_55_R0_data),
    .R0_en(mem_0_55_R0_en)
  );
  split_mem_ext mem_0_56 (
    .W0_addr(mem_0_56_W0_addr),
    .W0_clk(mem_0_56_W0_clk),
    .W0_data(mem_0_56_W0_data),
    .W0_en(mem_0_56_W0_en),
    .W0_mask(mem_0_56_W0_mask),
    .R0_addr(mem_0_56_R0_addr),
    .R0_clk(mem_0_56_R0_clk),
    .R0_data(mem_0_56_R0_data),
    .R0_en(mem_0_56_R0_en)
  );
  split_mem_ext mem_0_57 (
    .W0_addr(mem_0_57_W0_addr),
    .W0_clk(mem_0_57_W0_clk),
    .W0_data(mem_0_57_W0_data),
    .W0_en(mem_0_57_W0_en),
    .W0_mask(mem_0_57_W0_mask),
    .R0_addr(mem_0_57_R0_addr),
    .R0_clk(mem_0_57_R0_clk),
    .R0_data(mem_0_57_R0_data),
    .R0_en(mem_0_57_R0_en)
  );
  split_mem_ext mem_0_58 (
    .W0_addr(mem_0_58_W0_addr),
    .W0_clk(mem_0_58_W0_clk),
    .W0_data(mem_0_58_W0_data),
    .W0_en(mem_0_58_W0_en),
    .W0_mask(mem_0_58_W0_mask),
    .R0_addr(mem_0_58_R0_addr),
    .R0_clk(mem_0_58_R0_clk),
    .R0_data(mem_0_58_R0_data),
    .R0_en(mem_0_58_R0_en)
  );
  split_mem_ext mem_0_59 (
    .W0_addr(mem_0_59_W0_addr),
    .W0_clk(mem_0_59_W0_clk),
    .W0_data(mem_0_59_W0_data),
    .W0_en(mem_0_59_W0_en),
    .W0_mask(mem_0_59_W0_mask),
    .R0_addr(mem_0_59_R0_addr),
    .R0_clk(mem_0_59_R0_clk),
    .R0_data(mem_0_59_R0_data),
    .R0_en(mem_0_59_R0_en)
  );
  split_mem_ext mem_0_60 (
    .W0_addr(mem_0_60_W0_addr),
    .W0_clk(mem_0_60_W0_clk),
    .W0_data(mem_0_60_W0_data),
    .W0_en(mem_0_60_W0_en),
    .W0_mask(mem_0_60_W0_mask),
    .R0_addr(mem_0_60_R0_addr),
    .R0_clk(mem_0_60_R0_clk),
    .R0_data(mem_0_60_R0_data),
    .R0_en(mem_0_60_R0_en)
  );
  split_mem_ext mem_0_61 (
    .W0_addr(mem_0_61_W0_addr),
    .W0_clk(mem_0_61_W0_clk),
    .W0_data(mem_0_61_W0_data),
    .W0_en(mem_0_61_W0_en),
    .W0_mask(mem_0_61_W0_mask),
    .R0_addr(mem_0_61_R0_addr),
    .R0_clk(mem_0_61_R0_clk),
    .R0_data(mem_0_61_R0_data),
    .R0_en(mem_0_61_R0_en)
  );
  split_mem_ext mem_0_62 (
    .W0_addr(mem_0_62_W0_addr),
    .W0_clk(mem_0_62_W0_clk),
    .W0_data(mem_0_62_W0_data),
    .W0_en(mem_0_62_W0_en),
    .W0_mask(mem_0_62_W0_mask),
    .R0_addr(mem_0_62_R0_addr),
    .R0_clk(mem_0_62_R0_clk),
    .R0_data(mem_0_62_R0_data),
    .R0_en(mem_0_62_R0_en)
  );
  split_mem_ext mem_0_63 (
    .W0_addr(mem_0_63_W0_addr),
    .W0_clk(mem_0_63_W0_clk),
    .W0_data(mem_0_63_W0_data),
    .W0_en(mem_0_63_W0_en),
    .W0_mask(mem_0_63_W0_mask),
    .R0_addr(mem_0_63_R0_addr),
    .R0_clk(mem_0_63_R0_clk),
    .R0_data(mem_0_63_R0_data),
    .R0_en(mem_0_63_R0_en)
  );
  assign R0_data = {R0_data_0_63,_GEN_61};
  assign mem_0_0_W0_addr = W0_addr;
  assign mem_0_0_W0_clk = W0_clk;
  assign mem_0_0_W0_data = W0_data[7:0];
  assign mem_0_0_W0_en = W0_en;
  assign mem_0_0_W0_mask = W0_mask[0];
  assign mem_0_0_R0_addr = R0_addr;
  assign mem_0_0_R0_clk = R0_clk;
  assign mem_0_0_R0_en = R0_en;
  assign mem_0_1_W0_addr = W0_addr;
  assign mem_0_1_W0_clk = W0_clk;
  assign mem_0_1_W0_data = W0_data[15:8];
  assign mem_0_1_W0_en = W0_en;
  assign mem_0_1_W0_mask = W0_mask[1];
  assign mem_0_1_R0_addr = R0_addr;
  assign mem_0_1_R0_clk = R0_clk;
  assign mem_0_1_R0_en = R0_en;
  assign mem_0_2_W0_addr = W0_addr;
  assign mem_0_2_W0_clk = W0_clk;
  assign mem_0_2_W0_data = W0_data[23:16];
  assign mem_0_2_W0_en = W0_en;
  assign mem_0_2_W0_mask = W0_mask[2];
  assign mem_0_2_R0_addr = R0_addr;
  assign mem_0_2_R0_clk = R0_clk;
  assign mem_0_2_R0_en = R0_en;
  assign mem_0_3_W0_addr = W0_addr;
  assign mem_0_3_W0_clk = W0_clk;
  assign mem_0_3_W0_data = W0_data[31:24];
  assign mem_0_3_W0_en = W0_en;
  assign mem_0_3_W0_mask = W0_mask[3];
  assign mem_0_3_R0_addr = R0_addr;
  assign mem_0_3_R0_clk = R0_clk;
  assign mem_0_3_R0_en = R0_en;
  assign mem_0_4_W0_addr = W0_addr;
  assign mem_0_4_W0_clk = W0_clk;
  assign mem_0_4_W0_data = W0_data[39:32];
  assign mem_0_4_W0_en = W0_en;
  assign mem_0_4_W0_mask = W0_mask[4];
  assign mem_0_4_R0_addr = R0_addr;
  assign mem_0_4_R0_clk = R0_clk;
  assign mem_0_4_R0_en = R0_en;
  assign mem_0_5_W0_addr = W0_addr;
  assign mem_0_5_W0_clk = W0_clk;
  assign mem_0_5_W0_data = W0_data[47:40];
  assign mem_0_5_W0_en = W0_en;
  assign mem_0_5_W0_mask = W0_mask[5];
  assign mem_0_5_R0_addr = R0_addr;
  assign mem_0_5_R0_clk = R0_clk;
  assign mem_0_5_R0_en = R0_en;
  assign mem_0_6_W0_addr = W0_addr;
  assign mem_0_6_W0_clk = W0_clk;
  assign mem_0_6_W0_data = W0_data[55:48];
  assign mem_0_6_W0_en = W0_en;
  assign mem_0_6_W0_mask = W0_mask[6];
  assign mem_0_6_R0_addr = R0_addr;
  assign mem_0_6_R0_clk = R0_clk;
  assign mem_0_6_R0_en = R0_en;
  assign mem_0_7_W0_addr = W0_addr;
  assign mem_0_7_W0_clk = W0_clk;
  assign mem_0_7_W0_data = W0_data[63:56];
  assign mem_0_7_W0_en = W0_en;
  assign mem_0_7_W0_mask = W0_mask[7];
  assign mem_0_7_R0_addr = R0_addr;
  assign mem_0_7_R0_clk = R0_clk;
  assign mem_0_7_R0_en = R0_en;
  assign mem_0_8_W0_addr = W0_addr;
  assign mem_0_8_W0_clk = W0_clk;
  assign mem_0_8_W0_data = W0_data[71:64];
  assign mem_0_8_W0_en = W0_en;
  assign mem_0_8_W0_mask = W0_mask[8];
  assign mem_0_8_R0_addr = R0_addr;
  assign mem_0_8_R0_clk = R0_clk;
  assign mem_0_8_R0_en = R0_en;
  assign mem_0_9_W0_addr = W0_addr;
  assign mem_0_9_W0_clk = W0_clk;
  assign mem_0_9_W0_data = W0_data[79:72];
  assign mem_0_9_W0_en = W0_en;
  assign mem_0_9_W0_mask = W0_mask[9];
  assign mem_0_9_R0_addr = R0_addr;
  assign mem_0_9_R0_clk = R0_clk;
  assign mem_0_9_R0_en = R0_en;
  assign mem_0_10_W0_addr = W0_addr;
  assign mem_0_10_W0_clk = W0_clk;
  assign mem_0_10_W0_data = W0_data[87:80];
  assign mem_0_10_W0_en = W0_en;
  assign mem_0_10_W0_mask = W0_mask[10];
  assign mem_0_10_R0_addr = R0_addr;
  assign mem_0_10_R0_clk = R0_clk;
  assign mem_0_10_R0_en = R0_en;
  assign mem_0_11_W0_addr = W0_addr;
  assign mem_0_11_W0_clk = W0_clk;
  assign mem_0_11_W0_data = W0_data[95:88];
  assign mem_0_11_W0_en = W0_en;
  assign mem_0_11_W0_mask = W0_mask[11];
  assign mem_0_11_R0_addr = R0_addr;
  assign mem_0_11_R0_clk = R0_clk;
  assign mem_0_11_R0_en = R0_en;
  assign mem_0_12_W0_addr = W0_addr;
  assign mem_0_12_W0_clk = W0_clk;
  assign mem_0_12_W0_data = W0_data[103:96];
  assign mem_0_12_W0_en = W0_en;
  assign mem_0_12_W0_mask = W0_mask[12];
  assign mem_0_12_R0_addr = R0_addr;
  assign mem_0_12_R0_clk = R0_clk;
  assign mem_0_12_R0_en = R0_en;
  assign mem_0_13_W0_addr = W0_addr;
  assign mem_0_13_W0_clk = W0_clk;
  assign mem_0_13_W0_data = W0_data[111:104];
  assign mem_0_13_W0_en = W0_en;
  assign mem_0_13_W0_mask = W0_mask[13];
  assign mem_0_13_R0_addr = R0_addr;
  assign mem_0_13_R0_clk = R0_clk;
  assign mem_0_13_R0_en = R0_en;
  assign mem_0_14_W0_addr = W0_addr;
  assign mem_0_14_W0_clk = W0_clk;
  assign mem_0_14_W0_data = W0_data[119:112];
  assign mem_0_14_W0_en = W0_en;
  assign mem_0_14_W0_mask = W0_mask[14];
  assign mem_0_14_R0_addr = R0_addr;
  assign mem_0_14_R0_clk = R0_clk;
  assign mem_0_14_R0_en = R0_en;
  assign mem_0_15_W0_addr = W0_addr;
  assign mem_0_15_W0_clk = W0_clk;
  assign mem_0_15_W0_data = W0_data[127:120];
  assign mem_0_15_W0_en = W0_en;
  assign mem_0_15_W0_mask = W0_mask[15];
  assign mem_0_15_R0_addr = R0_addr;
  assign mem_0_15_R0_clk = R0_clk;
  assign mem_0_15_R0_en = R0_en;
  assign mem_0_16_W0_addr = W0_addr;
  assign mem_0_16_W0_clk = W0_clk;
  assign mem_0_16_W0_data = W0_data[135:128];
  assign mem_0_16_W0_en = W0_en;
  assign mem_0_16_W0_mask = W0_mask[16];
  assign mem_0_16_R0_addr = R0_addr;
  assign mem_0_16_R0_clk = R0_clk;
  assign mem_0_16_R0_en = R0_en;
  assign mem_0_17_W0_addr = W0_addr;
  assign mem_0_17_W0_clk = W0_clk;
  assign mem_0_17_W0_data = W0_data[143:136];
  assign mem_0_17_W0_en = W0_en;
  assign mem_0_17_W0_mask = W0_mask[17];
  assign mem_0_17_R0_addr = R0_addr;
  assign mem_0_17_R0_clk = R0_clk;
  assign mem_0_17_R0_en = R0_en;
  assign mem_0_18_W0_addr = W0_addr;
  assign mem_0_18_W0_clk = W0_clk;
  assign mem_0_18_W0_data = W0_data[151:144];
  assign mem_0_18_W0_en = W0_en;
  assign mem_0_18_W0_mask = W0_mask[18];
  assign mem_0_18_R0_addr = R0_addr;
  assign mem_0_18_R0_clk = R0_clk;
  assign mem_0_18_R0_en = R0_en;
  assign mem_0_19_W0_addr = W0_addr;
  assign mem_0_19_W0_clk = W0_clk;
  assign mem_0_19_W0_data = W0_data[159:152];
  assign mem_0_19_W0_en = W0_en;
  assign mem_0_19_W0_mask = W0_mask[19];
  assign mem_0_19_R0_addr = R0_addr;
  assign mem_0_19_R0_clk = R0_clk;
  assign mem_0_19_R0_en = R0_en;
  assign mem_0_20_W0_addr = W0_addr;
  assign mem_0_20_W0_clk = W0_clk;
  assign mem_0_20_W0_data = W0_data[167:160];
  assign mem_0_20_W0_en = W0_en;
  assign mem_0_20_W0_mask = W0_mask[20];
  assign mem_0_20_R0_addr = R0_addr;
  assign mem_0_20_R0_clk = R0_clk;
  assign mem_0_20_R0_en = R0_en;
  assign mem_0_21_W0_addr = W0_addr;
  assign mem_0_21_W0_clk = W0_clk;
  assign mem_0_21_W0_data = W0_data[175:168];
  assign mem_0_21_W0_en = W0_en;
  assign mem_0_21_W0_mask = W0_mask[21];
  assign mem_0_21_R0_addr = R0_addr;
  assign mem_0_21_R0_clk = R0_clk;
  assign mem_0_21_R0_en = R0_en;
  assign mem_0_22_W0_addr = W0_addr;
  assign mem_0_22_W0_clk = W0_clk;
  assign mem_0_22_W0_data = W0_data[183:176];
  assign mem_0_22_W0_en = W0_en;
  assign mem_0_22_W0_mask = W0_mask[22];
  assign mem_0_22_R0_addr = R0_addr;
  assign mem_0_22_R0_clk = R0_clk;
  assign mem_0_22_R0_en = R0_en;
  assign mem_0_23_W0_addr = W0_addr;
  assign mem_0_23_W0_clk = W0_clk;
  assign mem_0_23_W0_data = W0_data[191:184];
  assign mem_0_23_W0_en = W0_en;
  assign mem_0_23_W0_mask = W0_mask[23];
  assign mem_0_23_R0_addr = R0_addr;
  assign mem_0_23_R0_clk = R0_clk;
  assign mem_0_23_R0_en = R0_en;
  assign mem_0_24_W0_addr = W0_addr;
  assign mem_0_24_W0_clk = W0_clk;
  assign mem_0_24_W0_data = W0_data[199:192];
  assign mem_0_24_W0_en = W0_en;
  assign mem_0_24_W0_mask = W0_mask[24];
  assign mem_0_24_R0_addr = R0_addr;
  assign mem_0_24_R0_clk = R0_clk;
  assign mem_0_24_R0_en = R0_en;
  assign mem_0_25_W0_addr = W0_addr;
  assign mem_0_25_W0_clk = W0_clk;
  assign mem_0_25_W0_data = W0_data[207:200];
  assign mem_0_25_W0_en = W0_en;
  assign mem_0_25_W0_mask = W0_mask[25];
  assign mem_0_25_R0_addr = R0_addr;
  assign mem_0_25_R0_clk = R0_clk;
  assign mem_0_25_R0_en = R0_en;
  assign mem_0_26_W0_addr = W0_addr;
  assign mem_0_26_W0_clk = W0_clk;
  assign mem_0_26_W0_data = W0_data[215:208];
  assign mem_0_26_W0_en = W0_en;
  assign mem_0_26_W0_mask = W0_mask[26];
  assign mem_0_26_R0_addr = R0_addr;
  assign mem_0_26_R0_clk = R0_clk;
  assign mem_0_26_R0_en = R0_en;
  assign mem_0_27_W0_addr = W0_addr;
  assign mem_0_27_W0_clk = W0_clk;
  assign mem_0_27_W0_data = W0_data[223:216];
  assign mem_0_27_W0_en = W0_en;
  assign mem_0_27_W0_mask = W0_mask[27];
  assign mem_0_27_R0_addr = R0_addr;
  assign mem_0_27_R0_clk = R0_clk;
  assign mem_0_27_R0_en = R0_en;
  assign mem_0_28_W0_addr = W0_addr;
  assign mem_0_28_W0_clk = W0_clk;
  assign mem_0_28_W0_data = W0_data[231:224];
  assign mem_0_28_W0_en = W0_en;
  assign mem_0_28_W0_mask = W0_mask[28];
  assign mem_0_28_R0_addr = R0_addr;
  assign mem_0_28_R0_clk = R0_clk;
  assign mem_0_28_R0_en = R0_en;
  assign mem_0_29_W0_addr = W0_addr;
  assign mem_0_29_W0_clk = W0_clk;
  assign mem_0_29_W0_data = W0_data[239:232];
  assign mem_0_29_W0_en = W0_en;
  assign mem_0_29_W0_mask = W0_mask[29];
  assign mem_0_29_R0_addr = R0_addr;
  assign mem_0_29_R0_clk = R0_clk;
  assign mem_0_29_R0_en = R0_en;
  assign mem_0_30_W0_addr = W0_addr;
  assign mem_0_30_W0_clk = W0_clk;
  assign mem_0_30_W0_data = W0_data[247:240];
  assign mem_0_30_W0_en = W0_en;
  assign mem_0_30_W0_mask = W0_mask[30];
  assign mem_0_30_R0_addr = R0_addr;
  assign mem_0_30_R0_clk = R0_clk;
  assign mem_0_30_R0_en = R0_en;
  assign mem_0_31_W0_addr = W0_addr;
  assign mem_0_31_W0_clk = W0_clk;
  assign mem_0_31_W0_data = W0_data[255:248];
  assign mem_0_31_W0_en = W0_en;
  assign mem_0_31_W0_mask = W0_mask[31];
  assign mem_0_31_R0_addr = R0_addr;
  assign mem_0_31_R0_clk = R0_clk;
  assign mem_0_31_R0_en = R0_en;
  assign mem_0_32_W0_addr = W0_addr;
  assign mem_0_32_W0_clk = W0_clk;
  assign mem_0_32_W0_data = W0_data[263:256];
  assign mem_0_32_W0_en = W0_en;
  assign mem_0_32_W0_mask = W0_mask[32];
  assign mem_0_32_R0_addr = R0_addr;
  assign mem_0_32_R0_clk = R0_clk;
  assign mem_0_32_R0_en = R0_en;
  assign mem_0_33_W0_addr = W0_addr;
  assign mem_0_33_W0_clk = W0_clk;
  assign mem_0_33_W0_data = W0_data[271:264];
  assign mem_0_33_W0_en = W0_en;
  assign mem_0_33_W0_mask = W0_mask[33];
  assign mem_0_33_R0_addr = R0_addr;
  assign mem_0_33_R0_clk = R0_clk;
  assign mem_0_33_R0_en = R0_en;
  assign mem_0_34_W0_addr = W0_addr;
  assign mem_0_34_W0_clk = W0_clk;
  assign mem_0_34_W0_data = W0_data[279:272];
  assign mem_0_34_W0_en = W0_en;
  assign mem_0_34_W0_mask = W0_mask[34];
  assign mem_0_34_R0_addr = R0_addr;
  assign mem_0_34_R0_clk = R0_clk;
  assign mem_0_34_R0_en = R0_en;
  assign mem_0_35_W0_addr = W0_addr;
  assign mem_0_35_W0_clk = W0_clk;
  assign mem_0_35_W0_data = W0_data[287:280];
  assign mem_0_35_W0_en = W0_en;
  assign mem_0_35_W0_mask = W0_mask[35];
  assign mem_0_35_R0_addr = R0_addr;
  assign mem_0_35_R0_clk = R0_clk;
  assign mem_0_35_R0_en = R0_en;
  assign mem_0_36_W0_addr = W0_addr;
  assign mem_0_36_W0_clk = W0_clk;
  assign mem_0_36_W0_data = W0_data[295:288];
  assign mem_0_36_W0_en = W0_en;
  assign mem_0_36_W0_mask = W0_mask[36];
  assign mem_0_36_R0_addr = R0_addr;
  assign mem_0_36_R0_clk = R0_clk;
  assign mem_0_36_R0_en = R0_en;
  assign mem_0_37_W0_addr = W0_addr;
  assign mem_0_37_W0_clk = W0_clk;
  assign mem_0_37_W0_data = W0_data[303:296];
  assign mem_0_37_W0_en = W0_en;
  assign mem_0_37_W0_mask = W0_mask[37];
  assign mem_0_37_R0_addr = R0_addr;
  assign mem_0_37_R0_clk = R0_clk;
  assign mem_0_37_R0_en = R0_en;
  assign mem_0_38_W0_addr = W0_addr;
  assign mem_0_38_W0_clk = W0_clk;
  assign mem_0_38_W0_data = W0_data[311:304];
  assign mem_0_38_W0_en = W0_en;
  assign mem_0_38_W0_mask = W0_mask[38];
  assign mem_0_38_R0_addr = R0_addr;
  assign mem_0_38_R0_clk = R0_clk;
  assign mem_0_38_R0_en = R0_en;
  assign mem_0_39_W0_addr = W0_addr;
  assign mem_0_39_W0_clk = W0_clk;
  assign mem_0_39_W0_data = W0_data[319:312];
  assign mem_0_39_W0_en = W0_en;
  assign mem_0_39_W0_mask = W0_mask[39];
  assign mem_0_39_R0_addr = R0_addr;
  assign mem_0_39_R0_clk = R0_clk;
  assign mem_0_39_R0_en = R0_en;
  assign mem_0_40_W0_addr = W0_addr;
  assign mem_0_40_W0_clk = W0_clk;
  assign mem_0_40_W0_data = W0_data[327:320];
  assign mem_0_40_W0_en = W0_en;
  assign mem_0_40_W0_mask = W0_mask[40];
  assign mem_0_40_R0_addr = R0_addr;
  assign mem_0_40_R0_clk = R0_clk;
  assign mem_0_40_R0_en = R0_en;
  assign mem_0_41_W0_addr = W0_addr;
  assign mem_0_41_W0_clk = W0_clk;
  assign mem_0_41_W0_data = W0_data[335:328];
  assign mem_0_41_W0_en = W0_en;
  assign mem_0_41_W0_mask = W0_mask[41];
  assign mem_0_41_R0_addr = R0_addr;
  assign mem_0_41_R0_clk = R0_clk;
  assign mem_0_41_R0_en = R0_en;
  assign mem_0_42_W0_addr = W0_addr;
  assign mem_0_42_W0_clk = W0_clk;
  assign mem_0_42_W0_data = W0_data[343:336];
  assign mem_0_42_W0_en = W0_en;
  assign mem_0_42_W0_mask = W0_mask[42];
  assign mem_0_42_R0_addr = R0_addr;
  assign mem_0_42_R0_clk = R0_clk;
  assign mem_0_42_R0_en = R0_en;
  assign mem_0_43_W0_addr = W0_addr;
  assign mem_0_43_W0_clk = W0_clk;
  assign mem_0_43_W0_data = W0_data[351:344];
  assign mem_0_43_W0_en = W0_en;
  assign mem_0_43_W0_mask = W0_mask[43];
  assign mem_0_43_R0_addr = R0_addr;
  assign mem_0_43_R0_clk = R0_clk;
  assign mem_0_43_R0_en = R0_en;
  assign mem_0_44_W0_addr = W0_addr;
  assign mem_0_44_W0_clk = W0_clk;
  assign mem_0_44_W0_data = W0_data[359:352];
  assign mem_0_44_W0_en = W0_en;
  assign mem_0_44_W0_mask = W0_mask[44];
  assign mem_0_44_R0_addr = R0_addr;
  assign mem_0_44_R0_clk = R0_clk;
  assign mem_0_44_R0_en = R0_en;
  assign mem_0_45_W0_addr = W0_addr;
  assign mem_0_45_W0_clk = W0_clk;
  assign mem_0_45_W0_data = W0_data[367:360];
  assign mem_0_45_W0_en = W0_en;
  assign mem_0_45_W0_mask = W0_mask[45];
  assign mem_0_45_R0_addr = R0_addr;
  assign mem_0_45_R0_clk = R0_clk;
  assign mem_0_45_R0_en = R0_en;
  assign mem_0_46_W0_addr = W0_addr;
  assign mem_0_46_W0_clk = W0_clk;
  assign mem_0_46_W0_data = W0_data[375:368];
  assign mem_0_46_W0_en = W0_en;
  assign mem_0_46_W0_mask = W0_mask[46];
  assign mem_0_46_R0_addr = R0_addr;
  assign mem_0_46_R0_clk = R0_clk;
  assign mem_0_46_R0_en = R0_en;
  assign mem_0_47_W0_addr = W0_addr;
  assign mem_0_47_W0_clk = W0_clk;
  assign mem_0_47_W0_data = W0_data[383:376];
  assign mem_0_47_W0_en = W0_en;
  assign mem_0_47_W0_mask = W0_mask[47];
  assign mem_0_47_R0_addr = R0_addr;
  assign mem_0_47_R0_clk = R0_clk;
  assign mem_0_47_R0_en = R0_en;
  assign mem_0_48_W0_addr = W0_addr;
  assign mem_0_48_W0_clk = W0_clk;
  assign mem_0_48_W0_data = W0_data[391:384];
  assign mem_0_48_W0_en = W0_en;
  assign mem_0_48_W0_mask = W0_mask[48];
  assign mem_0_48_R0_addr = R0_addr;
  assign mem_0_48_R0_clk = R0_clk;
  assign mem_0_48_R0_en = R0_en;
  assign mem_0_49_W0_addr = W0_addr;
  assign mem_0_49_W0_clk = W0_clk;
  assign mem_0_49_W0_data = W0_data[399:392];
  assign mem_0_49_W0_en = W0_en;
  assign mem_0_49_W0_mask = W0_mask[49];
  assign mem_0_49_R0_addr = R0_addr;
  assign mem_0_49_R0_clk = R0_clk;
  assign mem_0_49_R0_en = R0_en;
  assign mem_0_50_W0_addr = W0_addr;
  assign mem_0_50_W0_clk = W0_clk;
  assign mem_0_50_W0_data = W0_data[407:400];
  assign mem_0_50_W0_en = W0_en;
  assign mem_0_50_W0_mask = W0_mask[50];
  assign mem_0_50_R0_addr = R0_addr;
  assign mem_0_50_R0_clk = R0_clk;
  assign mem_0_50_R0_en = R0_en;
  assign mem_0_51_W0_addr = W0_addr;
  assign mem_0_51_W0_clk = W0_clk;
  assign mem_0_51_W0_data = W0_data[415:408];
  assign mem_0_51_W0_en = W0_en;
  assign mem_0_51_W0_mask = W0_mask[51];
  assign mem_0_51_R0_addr = R0_addr;
  assign mem_0_51_R0_clk = R0_clk;
  assign mem_0_51_R0_en = R0_en;
  assign mem_0_52_W0_addr = W0_addr;
  assign mem_0_52_W0_clk = W0_clk;
  assign mem_0_52_W0_data = W0_data[423:416];
  assign mem_0_52_W0_en = W0_en;
  assign mem_0_52_W0_mask = W0_mask[52];
  assign mem_0_52_R0_addr = R0_addr;
  assign mem_0_52_R0_clk = R0_clk;
  assign mem_0_52_R0_en = R0_en;
  assign mem_0_53_W0_addr = W0_addr;
  assign mem_0_53_W0_clk = W0_clk;
  assign mem_0_53_W0_data = W0_data[431:424];
  assign mem_0_53_W0_en = W0_en;
  assign mem_0_53_W0_mask = W0_mask[53];
  assign mem_0_53_R0_addr = R0_addr;
  assign mem_0_53_R0_clk = R0_clk;
  assign mem_0_53_R0_en = R0_en;
  assign mem_0_54_W0_addr = W0_addr;
  assign mem_0_54_W0_clk = W0_clk;
  assign mem_0_54_W0_data = W0_data[439:432];
  assign mem_0_54_W0_en = W0_en;
  assign mem_0_54_W0_mask = W0_mask[54];
  assign mem_0_54_R0_addr = R0_addr;
  assign mem_0_54_R0_clk = R0_clk;
  assign mem_0_54_R0_en = R0_en;
  assign mem_0_55_W0_addr = W0_addr;
  assign mem_0_55_W0_clk = W0_clk;
  assign mem_0_55_W0_data = W0_data[447:440];
  assign mem_0_55_W0_en = W0_en;
  assign mem_0_55_W0_mask = W0_mask[55];
  assign mem_0_55_R0_addr = R0_addr;
  assign mem_0_55_R0_clk = R0_clk;
  assign mem_0_55_R0_en = R0_en;
  assign mem_0_56_W0_addr = W0_addr;
  assign mem_0_56_W0_clk = W0_clk;
  assign mem_0_56_W0_data = W0_data[455:448];
  assign mem_0_56_W0_en = W0_en;
  assign mem_0_56_W0_mask = W0_mask[56];
  assign mem_0_56_R0_addr = R0_addr;
  assign mem_0_56_R0_clk = R0_clk;
  assign mem_0_56_R0_en = R0_en;
  assign mem_0_57_W0_addr = W0_addr;
  assign mem_0_57_W0_clk = W0_clk;
  assign mem_0_57_W0_data = W0_data[463:456];
  assign mem_0_57_W0_en = W0_en;
  assign mem_0_57_W0_mask = W0_mask[57];
  assign mem_0_57_R0_addr = R0_addr;
  assign mem_0_57_R0_clk = R0_clk;
  assign mem_0_57_R0_en = R0_en;
  assign mem_0_58_W0_addr = W0_addr;
  assign mem_0_58_W0_clk = W0_clk;
  assign mem_0_58_W0_data = W0_data[471:464];
  assign mem_0_58_W0_en = W0_en;
  assign mem_0_58_W0_mask = W0_mask[58];
  assign mem_0_58_R0_addr = R0_addr;
  assign mem_0_58_R0_clk = R0_clk;
  assign mem_0_58_R0_en = R0_en;
  assign mem_0_59_W0_addr = W0_addr;
  assign mem_0_59_W0_clk = W0_clk;
  assign mem_0_59_W0_data = W0_data[479:472];
  assign mem_0_59_W0_en = W0_en;
  assign mem_0_59_W0_mask = W0_mask[59];
  assign mem_0_59_R0_addr = R0_addr;
  assign mem_0_59_R0_clk = R0_clk;
  assign mem_0_59_R0_en = R0_en;
  assign mem_0_60_W0_addr = W0_addr;
  assign mem_0_60_W0_clk = W0_clk;
  assign mem_0_60_W0_data = W0_data[487:480];
  assign mem_0_60_W0_en = W0_en;
  assign mem_0_60_W0_mask = W0_mask[60];
  assign mem_0_60_R0_addr = R0_addr;
  assign mem_0_60_R0_clk = R0_clk;
  assign mem_0_60_R0_en = R0_en;
  assign mem_0_61_W0_addr = W0_addr;
  assign mem_0_61_W0_clk = W0_clk;
  assign mem_0_61_W0_data = W0_data[495:488];
  assign mem_0_61_W0_en = W0_en;
  assign mem_0_61_W0_mask = W0_mask[61];
  assign mem_0_61_R0_addr = R0_addr;
  assign mem_0_61_R0_clk = R0_clk;
  assign mem_0_61_R0_en = R0_en;
  assign mem_0_62_W0_addr = W0_addr;
  assign mem_0_62_W0_clk = W0_clk;
  assign mem_0_62_W0_data = W0_data[503:496];
  assign mem_0_62_W0_en = W0_en;
  assign mem_0_62_W0_mask = W0_mask[62];
  assign mem_0_62_R0_addr = R0_addr;
  assign mem_0_62_R0_clk = R0_clk;
  assign mem_0_62_R0_en = R0_en;
  assign mem_0_63_W0_addr = W0_addr;
  assign mem_0_63_W0_clk = W0_clk;
  assign mem_0_63_W0_data = W0_data[511:504];
  assign mem_0_63_W0_en = W0_en;
  assign mem_0_63_W0_mask = W0_mask[63];
  assign mem_0_63_R0_addr = R0_addr;
  assign mem_0_63_R0_clk = R0_clk;
  assign mem_0_63_R0_en = R0_en;
endmodule
module mem_0_ext(
  input  [6:0]    W0_addr,
  input           W0_clk,
  input  [2047:0] W0_data,
  input           W0_en,
  input  [255:0]  W0_mask,
  input  [6:0]    R0_addr,
  input           R0_clk,
  output [2047:0] R0_data,
  input           R0_en
);
  wire [6:0] mem_0_0_W0_addr;
  wire  mem_0_0_W0_clk;
  wire [7:0] mem_0_0_W0_data;
  wire  mem_0_0_W0_en;
  wire  mem_0_0_W0_mask;
  wire [6:0] mem_0_0_R0_addr;
  wire  mem_0_0_R0_clk;
  wire [7:0] mem_0_0_R0_data;
  wire  mem_0_0_R0_en;
  wire [6:0] mem_0_1_W0_addr;
  wire  mem_0_1_W0_clk;
  wire [7:0] mem_0_1_W0_data;
  wire  mem_0_1_W0_en;
  wire  mem_0_1_W0_mask;
  wire [6:0] mem_0_1_R0_addr;
  wire  mem_0_1_R0_clk;
  wire [7:0] mem_0_1_R0_data;
  wire  mem_0_1_R0_en;
  wire [6:0] mem_0_2_W0_addr;
  wire  mem_0_2_W0_clk;
  wire [7:0] mem_0_2_W0_data;
  wire  mem_0_2_W0_en;
  wire  mem_0_2_W0_mask;
  wire [6:0] mem_0_2_R0_addr;
  wire  mem_0_2_R0_clk;
  wire [7:0] mem_0_2_R0_data;
  wire  mem_0_2_R0_en;
  wire [6:0] mem_0_3_W0_addr;
  wire  mem_0_3_W0_clk;
  wire [7:0] mem_0_3_W0_data;
  wire  mem_0_3_W0_en;
  wire  mem_0_3_W0_mask;
  wire [6:0] mem_0_3_R0_addr;
  wire  mem_0_3_R0_clk;
  wire [7:0] mem_0_3_R0_data;
  wire  mem_0_3_R0_en;
  wire [6:0] mem_0_4_W0_addr;
  wire  mem_0_4_W0_clk;
  wire [7:0] mem_0_4_W0_data;
  wire  mem_0_4_W0_en;
  wire  mem_0_4_W0_mask;
  wire [6:0] mem_0_4_R0_addr;
  wire  mem_0_4_R0_clk;
  wire [7:0] mem_0_4_R0_data;
  wire  mem_0_4_R0_en;
  wire [6:0] mem_0_5_W0_addr;
  wire  mem_0_5_W0_clk;
  wire [7:0] mem_0_5_W0_data;
  wire  mem_0_5_W0_en;
  wire  mem_0_5_W0_mask;
  wire [6:0] mem_0_5_R0_addr;
  wire  mem_0_5_R0_clk;
  wire [7:0] mem_0_5_R0_data;
  wire  mem_0_5_R0_en;
  wire [6:0] mem_0_6_W0_addr;
  wire  mem_0_6_W0_clk;
  wire [7:0] mem_0_6_W0_data;
  wire  mem_0_6_W0_en;
  wire  mem_0_6_W0_mask;
  wire [6:0] mem_0_6_R0_addr;
  wire  mem_0_6_R0_clk;
  wire [7:0] mem_0_6_R0_data;
  wire  mem_0_6_R0_en;
  wire [6:0] mem_0_7_W0_addr;
  wire  mem_0_7_W0_clk;
  wire [7:0] mem_0_7_W0_data;
  wire  mem_0_7_W0_en;
  wire  mem_0_7_W0_mask;
  wire [6:0] mem_0_7_R0_addr;
  wire  mem_0_7_R0_clk;
  wire [7:0] mem_0_7_R0_data;
  wire  mem_0_7_R0_en;
  wire [6:0] mem_0_8_W0_addr;
  wire  mem_0_8_W0_clk;
  wire [7:0] mem_0_8_W0_data;
  wire  mem_0_8_W0_en;
  wire  mem_0_8_W0_mask;
  wire [6:0] mem_0_8_R0_addr;
  wire  mem_0_8_R0_clk;
  wire [7:0] mem_0_8_R0_data;
  wire  mem_0_8_R0_en;
  wire [6:0] mem_0_9_W0_addr;
  wire  mem_0_9_W0_clk;
  wire [7:0] mem_0_9_W0_data;
  wire  mem_0_9_W0_en;
  wire  mem_0_9_W0_mask;
  wire [6:0] mem_0_9_R0_addr;
  wire  mem_0_9_R0_clk;
  wire [7:0] mem_0_9_R0_data;
  wire  mem_0_9_R0_en;
  wire [6:0] mem_0_10_W0_addr;
  wire  mem_0_10_W0_clk;
  wire [7:0] mem_0_10_W0_data;
  wire  mem_0_10_W0_en;
  wire  mem_0_10_W0_mask;
  wire [6:0] mem_0_10_R0_addr;
  wire  mem_0_10_R0_clk;
  wire [7:0] mem_0_10_R0_data;
  wire  mem_0_10_R0_en;
  wire [6:0] mem_0_11_W0_addr;
  wire  mem_0_11_W0_clk;
  wire [7:0] mem_0_11_W0_data;
  wire  mem_0_11_W0_en;
  wire  mem_0_11_W0_mask;
  wire [6:0] mem_0_11_R0_addr;
  wire  mem_0_11_R0_clk;
  wire [7:0] mem_0_11_R0_data;
  wire  mem_0_11_R0_en;
  wire [6:0] mem_0_12_W0_addr;
  wire  mem_0_12_W0_clk;
  wire [7:0] mem_0_12_W0_data;
  wire  mem_0_12_W0_en;
  wire  mem_0_12_W0_mask;
  wire [6:0] mem_0_12_R0_addr;
  wire  mem_0_12_R0_clk;
  wire [7:0] mem_0_12_R0_data;
  wire  mem_0_12_R0_en;
  wire [6:0] mem_0_13_W0_addr;
  wire  mem_0_13_W0_clk;
  wire [7:0] mem_0_13_W0_data;
  wire  mem_0_13_W0_en;
  wire  mem_0_13_W0_mask;
  wire [6:0] mem_0_13_R0_addr;
  wire  mem_0_13_R0_clk;
  wire [7:0] mem_0_13_R0_data;
  wire  mem_0_13_R0_en;
  wire [6:0] mem_0_14_W0_addr;
  wire  mem_0_14_W0_clk;
  wire [7:0] mem_0_14_W0_data;
  wire  mem_0_14_W0_en;
  wire  mem_0_14_W0_mask;
  wire [6:0] mem_0_14_R0_addr;
  wire  mem_0_14_R0_clk;
  wire [7:0] mem_0_14_R0_data;
  wire  mem_0_14_R0_en;
  wire [6:0] mem_0_15_W0_addr;
  wire  mem_0_15_W0_clk;
  wire [7:0] mem_0_15_W0_data;
  wire  mem_0_15_W0_en;
  wire  mem_0_15_W0_mask;
  wire [6:0] mem_0_15_R0_addr;
  wire  mem_0_15_R0_clk;
  wire [7:0] mem_0_15_R0_data;
  wire  mem_0_15_R0_en;
  wire [6:0] mem_0_16_W0_addr;
  wire  mem_0_16_W0_clk;
  wire [7:0] mem_0_16_W0_data;
  wire  mem_0_16_W0_en;
  wire  mem_0_16_W0_mask;
  wire [6:0] mem_0_16_R0_addr;
  wire  mem_0_16_R0_clk;
  wire [7:0] mem_0_16_R0_data;
  wire  mem_0_16_R0_en;
  wire [6:0] mem_0_17_W0_addr;
  wire  mem_0_17_W0_clk;
  wire [7:0] mem_0_17_W0_data;
  wire  mem_0_17_W0_en;
  wire  mem_0_17_W0_mask;
  wire [6:0] mem_0_17_R0_addr;
  wire  mem_0_17_R0_clk;
  wire [7:0] mem_0_17_R0_data;
  wire  mem_0_17_R0_en;
  wire [6:0] mem_0_18_W0_addr;
  wire  mem_0_18_W0_clk;
  wire [7:0] mem_0_18_W0_data;
  wire  mem_0_18_W0_en;
  wire  mem_0_18_W0_mask;
  wire [6:0] mem_0_18_R0_addr;
  wire  mem_0_18_R0_clk;
  wire [7:0] mem_0_18_R0_data;
  wire  mem_0_18_R0_en;
  wire [6:0] mem_0_19_W0_addr;
  wire  mem_0_19_W0_clk;
  wire [7:0] mem_0_19_W0_data;
  wire  mem_0_19_W0_en;
  wire  mem_0_19_W0_mask;
  wire [6:0] mem_0_19_R0_addr;
  wire  mem_0_19_R0_clk;
  wire [7:0] mem_0_19_R0_data;
  wire  mem_0_19_R0_en;
  wire [6:0] mem_0_20_W0_addr;
  wire  mem_0_20_W0_clk;
  wire [7:0] mem_0_20_W0_data;
  wire  mem_0_20_W0_en;
  wire  mem_0_20_W0_mask;
  wire [6:0] mem_0_20_R0_addr;
  wire  mem_0_20_R0_clk;
  wire [7:0] mem_0_20_R0_data;
  wire  mem_0_20_R0_en;
  wire [6:0] mem_0_21_W0_addr;
  wire  mem_0_21_W0_clk;
  wire [7:0] mem_0_21_W0_data;
  wire  mem_0_21_W0_en;
  wire  mem_0_21_W0_mask;
  wire [6:0] mem_0_21_R0_addr;
  wire  mem_0_21_R0_clk;
  wire [7:0] mem_0_21_R0_data;
  wire  mem_0_21_R0_en;
  wire [6:0] mem_0_22_W0_addr;
  wire  mem_0_22_W0_clk;
  wire [7:0] mem_0_22_W0_data;
  wire  mem_0_22_W0_en;
  wire  mem_0_22_W0_mask;
  wire [6:0] mem_0_22_R0_addr;
  wire  mem_0_22_R0_clk;
  wire [7:0] mem_0_22_R0_data;
  wire  mem_0_22_R0_en;
  wire [6:0] mem_0_23_W0_addr;
  wire  mem_0_23_W0_clk;
  wire [7:0] mem_0_23_W0_data;
  wire  mem_0_23_W0_en;
  wire  mem_0_23_W0_mask;
  wire [6:0] mem_0_23_R0_addr;
  wire  mem_0_23_R0_clk;
  wire [7:0] mem_0_23_R0_data;
  wire  mem_0_23_R0_en;
  wire [6:0] mem_0_24_W0_addr;
  wire  mem_0_24_W0_clk;
  wire [7:0] mem_0_24_W0_data;
  wire  mem_0_24_W0_en;
  wire  mem_0_24_W0_mask;
  wire [6:0] mem_0_24_R0_addr;
  wire  mem_0_24_R0_clk;
  wire [7:0] mem_0_24_R0_data;
  wire  mem_0_24_R0_en;
  wire [6:0] mem_0_25_W0_addr;
  wire  mem_0_25_W0_clk;
  wire [7:0] mem_0_25_W0_data;
  wire  mem_0_25_W0_en;
  wire  mem_0_25_W0_mask;
  wire [6:0] mem_0_25_R0_addr;
  wire  mem_0_25_R0_clk;
  wire [7:0] mem_0_25_R0_data;
  wire  mem_0_25_R0_en;
  wire [6:0] mem_0_26_W0_addr;
  wire  mem_0_26_W0_clk;
  wire [7:0] mem_0_26_W0_data;
  wire  mem_0_26_W0_en;
  wire  mem_0_26_W0_mask;
  wire [6:0] mem_0_26_R0_addr;
  wire  mem_0_26_R0_clk;
  wire [7:0] mem_0_26_R0_data;
  wire  mem_0_26_R0_en;
  wire [6:0] mem_0_27_W0_addr;
  wire  mem_0_27_W0_clk;
  wire [7:0] mem_0_27_W0_data;
  wire  mem_0_27_W0_en;
  wire  mem_0_27_W0_mask;
  wire [6:0] mem_0_27_R0_addr;
  wire  mem_0_27_R0_clk;
  wire [7:0] mem_0_27_R0_data;
  wire  mem_0_27_R0_en;
  wire [6:0] mem_0_28_W0_addr;
  wire  mem_0_28_W0_clk;
  wire [7:0] mem_0_28_W0_data;
  wire  mem_0_28_W0_en;
  wire  mem_0_28_W0_mask;
  wire [6:0] mem_0_28_R0_addr;
  wire  mem_0_28_R0_clk;
  wire [7:0] mem_0_28_R0_data;
  wire  mem_0_28_R0_en;
  wire [6:0] mem_0_29_W0_addr;
  wire  mem_0_29_W0_clk;
  wire [7:0] mem_0_29_W0_data;
  wire  mem_0_29_W0_en;
  wire  mem_0_29_W0_mask;
  wire [6:0] mem_0_29_R0_addr;
  wire  mem_0_29_R0_clk;
  wire [7:0] mem_0_29_R0_data;
  wire  mem_0_29_R0_en;
  wire [6:0] mem_0_30_W0_addr;
  wire  mem_0_30_W0_clk;
  wire [7:0] mem_0_30_W0_data;
  wire  mem_0_30_W0_en;
  wire  mem_0_30_W0_mask;
  wire [6:0] mem_0_30_R0_addr;
  wire  mem_0_30_R0_clk;
  wire [7:0] mem_0_30_R0_data;
  wire  mem_0_30_R0_en;
  wire [6:0] mem_0_31_W0_addr;
  wire  mem_0_31_W0_clk;
  wire [7:0] mem_0_31_W0_data;
  wire  mem_0_31_W0_en;
  wire  mem_0_31_W0_mask;
  wire [6:0] mem_0_31_R0_addr;
  wire  mem_0_31_R0_clk;
  wire [7:0] mem_0_31_R0_data;
  wire  mem_0_31_R0_en;
  wire [6:0] mem_0_32_W0_addr;
  wire  mem_0_32_W0_clk;
  wire [7:0] mem_0_32_W0_data;
  wire  mem_0_32_W0_en;
  wire  mem_0_32_W0_mask;
  wire [6:0] mem_0_32_R0_addr;
  wire  mem_0_32_R0_clk;
  wire [7:0] mem_0_32_R0_data;
  wire  mem_0_32_R0_en;
  wire [6:0] mem_0_33_W0_addr;
  wire  mem_0_33_W0_clk;
  wire [7:0] mem_0_33_W0_data;
  wire  mem_0_33_W0_en;
  wire  mem_0_33_W0_mask;
  wire [6:0] mem_0_33_R0_addr;
  wire  mem_0_33_R0_clk;
  wire [7:0] mem_0_33_R0_data;
  wire  mem_0_33_R0_en;
  wire [6:0] mem_0_34_W0_addr;
  wire  mem_0_34_W0_clk;
  wire [7:0] mem_0_34_W0_data;
  wire  mem_0_34_W0_en;
  wire  mem_0_34_W0_mask;
  wire [6:0] mem_0_34_R0_addr;
  wire  mem_0_34_R0_clk;
  wire [7:0] mem_0_34_R0_data;
  wire  mem_0_34_R0_en;
  wire [6:0] mem_0_35_W0_addr;
  wire  mem_0_35_W0_clk;
  wire [7:0] mem_0_35_W0_data;
  wire  mem_0_35_W0_en;
  wire  mem_0_35_W0_mask;
  wire [6:0] mem_0_35_R0_addr;
  wire  mem_0_35_R0_clk;
  wire [7:0] mem_0_35_R0_data;
  wire  mem_0_35_R0_en;
  wire [6:0] mem_0_36_W0_addr;
  wire  mem_0_36_W0_clk;
  wire [7:0] mem_0_36_W0_data;
  wire  mem_0_36_W0_en;
  wire  mem_0_36_W0_mask;
  wire [6:0] mem_0_36_R0_addr;
  wire  mem_0_36_R0_clk;
  wire [7:0] mem_0_36_R0_data;
  wire  mem_0_36_R0_en;
  wire [6:0] mem_0_37_W0_addr;
  wire  mem_0_37_W0_clk;
  wire [7:0] mem_0_37_W0_data;
  wire  mem_0_37_W0_en;
  wire  mem_0_37_W0_mask;
  wire [6:0] mem_0_37_R0_addr;
  wire  mem_0_37_R0_clk;
  wire [7:0] mem_0_37_R0_data;
  wire  mem_0_37_R0_en;
  wire [6:0] mem_0_38_W0_addr;
  wire  mem_0_38_W0_clk;
  wire [7:0] mem_0_38_W0_data;
  wire  mem_0_38_W0_en;
  wire  mem_0_38_W0_mask;
  wire [6:0] mem_0_38_R0_addr;
  wire  mem_0_38_R0_clk;
  wire [7:0] mem_0_38_R0_data;
  wire  mem_0_38_R0_en;
  wire [6:0] mem_0_39_W0_addr;
  wire  mem_0_39_W0_clk;
  wire [7:0] mem_0_39_W0_data;
  wire  mem_0_39_W0_en;
  wire  mem_0_39_W0_mask;
  wire [6:0] mem_0_39_R0_addr;
  wire  mem_0_39_R0_clk;
  wire [7:0] mem_0_39_R0_data;
  wire  mem_0_39_R0_en;
  wire [6:0] mem_0_40_W0_addr;
  wire  mem_0_40_W0_clk;
  wire [7:0] mem_0_40_W0_data;
  wire  mem_0_40_W0_en;
  wire  mem_0_40_W0_mask;
  wire [6:0] mem_0_40_R0_addr;
  wire  mem_0_40_R0_clk;
  wire [7:0] mem_0_40_R0_data;
  wire  mem_0_40_R0_en;
  wire [6:0] mem_0_41_W0_addr;
  wire  mem_0_41_W0_clk;
  wire [7:0] mem_0_41_W0_data;
  wire  mem_0_41_W0_en;
  wire  mem_0_41_W0_mask;
  wire [6:0] mem_0_41_R0_addr;
  wire  mem_0_41_R0_clk;
  wire [7:0] mem_0_41_R0_data;
  wire  mem_0_41_R0_en;
  wire [6:0] mem_0_42_W0_addr;
  wire  mem_0_42_W0_clk;
  wire [7:0] mem_0_42_W0_data;
  wire  mem_0_42_W0_en;
  wire  mem_0_42_W0_mask;
  wire [6:0] mem_0_42_R0_addr;
  wire  mem_0_42_R0_clk;
  wire [7:0] mem_0_42_R0_data;
  wire  mem_0_42_R0_en;
  wire [6:0] mem_0_43_W0_addr;
  wire  mem_0_43_W0_clk;
  wire [7:0] mem_0_43_W0_data;
  wire  mem_0_43_W0_en;
  wire  mem_0_43_W0_mask;
  wire [6:0] mem_0_43_R0_addr;
  wire  mem_0_43_R0_clk;
  wire [7:0] mem_0_43_R0_data;
  wire  mem_0_43_R0_en;
  wire [6:0] mem_0_44_W0_addr;
  wire  mem_0_44_W0_clk;
  wire [7:0] mem_0_44_W0_data;
  wire  mem_0_44_W0_en;
  wire  mem_0_44_W0_mask;
  wire [6:0] mem_0_44_R0_addr;
  wire  mem_0_44_R0_clk;
  wire [7:0] mem_0_44_R0_data;
  wire  mem_0_44_R0_en;
  wire [6:0] mem_0_45_W0_addr;
  wire  mem_0_45_W0_clk;
  wire [7:0] mem_0_45_W0_data;
  wire  mem_0_45_W0_en;
  wire  mem_0_45_W0_mask;
  wire [6:0] mem_0_45_R0_addr;
  wire  mem_0_45_R0_clk;
  wire [7:0] mem_0_45_R0_data;
  wire  mem_0_45_R0_en;
  wire [6:0] mem_0_46_W0_addr;
  wire  mem_0_46_W0_clk;
  wire [7:0] mem_0_46_W0_data;
  wire  mem_0_46_W0_en;
  wire  mem_0_46_W0_mask;
  wire [6:0] mem_0_46_R0_addr;
  wire  mem_0_46_R0_clk;
  wire [7:0] mem_0_46_R0_data;
  wire  mem_0_46_R0_en;
  wire [6:0] mem_0_47_W0_addr;
  wire  mem_0_47_W0_clk;
  wire [7:0] mem_0_47_W0_data;
  wire  mem_0_47_W0_en;
  wire  mem_0_47_W0_mask;
  wire [6:0] mem_0_47_R0_addr;
  wire  mem_0_47_R0_clk;
  wire [7:0] mem_0_47_R0_data;
  wire  mem_0_47_R0_en;
  wire [6:0] mem_0_48_W0_addr;
  wire  mem_0_48_W0_clk;
  wire [7:0] mem_0_48_W0_data;
  wire  mem_0_48_W0_en;
  wire  mem_0_48_W0_mask;
  wire [6:0] mem_0_48_R0_addr;
  wire  mem_0_48_R0_clk;
  wire [7:0] mem_0_48_R0_data;
  wire  mem_0_48_R0_en;
  wire [6:0] mem_0_49_W0_addr;
  wire  mem_0_49_W0_clk;
  wire [7:0] mem_0_49_W0_data;
  wire  mem_0_49_W0_en;
  wire  mem_0_49_W0_mask;
  wire [6:0] mem_0_49_R0_addr;
  wire  mem_0_49_R0_clk;
  wire [7:0] mem_0_49_R0_data;
  wire  mem_0_49_R0_en;
  wire [6:0] mem_0_50_W0_addr;
  wire  mem_0_50_W0_clk;
  wire [7:0] mem_0_50_W0_data;
  wire  mem_0_50_W0_en;
  wire  mem_0_50_W0_mask;
  wire [6:0] mem_0_50_R0_addr;
  wire  mem_0_50_R0_clk;
  wire [7:0] mem_0_50_R0_data;
  wire  mem_0_50_R0_en;
  wire [6:0] mem_0_51_W0_addr;
  wire  mem_0_51_W0_clk;
  wire [7:0] mem_0_51_W0_data;
  wire  mem_0_51_W0_en;
  wire  mem_0_51_W0_mask;
  wire [6:0] mem_0_51_R0_addr;
  wire  mem_0_51_R0_clk;
  wire [7:0] mem_0_51_R0_data;
  wire  mem_0_51_R0_en;
  wire [6:0] mem_0_52_W0_addr;
  wire  mem_0_52_W0_clk;
  wire [7:0] mem_0_52_W0_data;
  wire  mem_0_52_W0_en;
  wire  mem_0_52_W0_mask;
  wire [6:0] mem_0_52_R0_addr;
  wire  mem_0_52_R0_clk;
  wire [7:0] mem_0_52_R0_data;
  wire  mem_0_52_R0_en;
  wire [6:0] mem_0_53_W0_addr;
  wire  mem_0_53_W0_clk;
  wire [7:0] mem_0_53_W0_data;
  wire  mem_0_53_W0_en;
  wire  mem_0_53_W0_mask;
  wire [6:0] mem_0_53_R0_addr;
  wire  mem_0_53_R0_clk;
  wire [7:0] mem_0_53_R0_data;
  wire  mem_0_53_R0_en;
  wire [6:0] mem_0_54_W0_addr;
  wire  mem_0_54_W0_clk;
  wire [7:0] mem_0_54_W0_data;
  wire  mem_0_54_W0_en;
  wire  mem_0_54_W0_mask;
  wire [6:0] mem_0_54_R0_addr;
  wire  mem_0_54_R0_clk;
  wire [7:0] mem_0_54_R0_data;
  wire  mem_0_54_R0_en;
  wire [6:0] mem_0_55_W0_addr;
  wire  mem_0_55_W0_clk;
  wire [7:0] mem_0_55_W0_data;
  wire  mem_0_55_W0_en;
  wire  mem_0_55_W0_mask;
  wire [6:0] mem_0_55_R0_addr;
  wire  mem_0_55_R0_clk;
  wire [7:0] mem_0_55_R0_data;
  wire  mem_0_55_R0_en;
  wire [6:0] mem_0_56_W0_addr;
  wire  mem_0_56_W0_clk;
  wire [7:0] mem_0_56_W0_data;
  wire  mem_0_56_W0_en;
  wire  mem_0_56_W0_mask;
  wire [6:0] mem_0_56_R0_addr;
  wire  mem_0_56_R0_clk;
  wire [7:0] mem_0_56_R0_data;
  wire  mem_0_56_R0_en;
  wire [6:0] mem_0_57_W0_addr;
  wire  mem_0_57_W0_clk;
  wire [7:0] mem_0_57_W0_data;
  wire  mem_0_57_W0_en;
  wire  mem_0_57_W0_mask;
  wire [6:0] mem_0_57_R0_addr;
  wire  mem_0_57_R0_clk;
  wire [7:0] mem_0_57_R0_data;
  wire  mem_0_57_R0_en;
  wire [6:0] mem_0_58_W0_addr;
  wire  mem_0_58_W0_clk;
  wire [7:0] mem_0_58_W0_data;
  wire  mem_0_58_W0_en;
  wire  mem_0_58_W0_mask;
  wire [6:0] mem_0_58_R0_addr;
  wire  mem_0_58_R0_clk;
  wire [7:0] mem_0_58_R0_data;
  wire  mem_0_58_R0_en;
  wire [6:0] mem_0_59_W0_addr;
  wire  mem_0_59_W0_clk;
  wire [7:0] mem_0_59_W0_data;
  wire  mem_0_59_W0_en;
  wire  mem_0_59_W0_mask;
  wire [6:0] mem_0_59_R0_addr;
  wire  mem_0_59_R0_clk;
  wire [7:0] mem_0_59_R0_data;
  wire  mem_0_59_R0_en;
  wire [6:0] mem_0_60_W0_addr;
  wire  mem_0_60_W0_clk;
  wire [7:0] mem_0_60_W0_data;
  wire  mem_0_60_W0_en;
  wire  mem_0_60_W0_mask;
  wire [6:0] mem_0_60_R0_addr;
  wire  mem_0_60_R0_clk;
  wire [7:0] mem_0_60_R0_data;
  wire  mem_0_60_R0_en;
  wire [6:0] mem_0_61_W0_addr;
  wire  mem_0_61_W0_clk;
  wire [7:0] mem_0_61_W0_data;
  wire  mem_0_61_W0_en;
  wire  mem_0_61_W0_mask;
  wire [6:0] mem_0_61_R0_addr;
  wire  mem_0_61_R0_clk;
  wire [7:0] mem_0_61_R0_data;
  wire  mem_0_61_R0_en;
  wire [6:0] mem_0_62_W0_addr;
  wire  mem_0_62_W0_clk;
  wire [7:0] mem_0_62_W0_data;
  wire  mem_0_62_W0_en;
  wire  mem_0_62_W0_mask;
  wire [6:0] mem_0_62_R0_addr;
  wire  mem_0_62_R0_clk;
  wire [7:0] mem_0_62_R0_data;
  wire  mem_0_62_R0_en;
  wire [6:0] mem_0_63_W0_addr;
  wire  mem_0_63_W0_clk;
  wire [7:0] mem_0_63_W0_data;
  wire  mem_0_63_W0_en;
  wire  mem_0_63_W0_mask;
  wire [6:0] mem_0_63_R0_addr;
  wire  mem_0_63_R0_clk;
  wire [7:0] mem_0_63_R0_data;
  wire  mem_0_63_R0_en;
  wire [6:0] mem_0_64_W0_addr;
  wire  mem_0_64_W0_clk;
  wire [7:0] mem_0_64_W0_data;
  wire  mem_0_64_W0_en;
  wire  mem_0_64_W0_mask;
  wire [6:0] mem_0_64_R0_addr;
  wire  mem_0_64_R0_clk;
  wire [7:0] mem_0_64_R0_data;
  wire  mem_0_64_R0_en;
  wire [6:0] mem_0_65_W0_addr;
  wire  mem_0_65_W0_clk;
  wire [7:0] mem_0_65_W0_data;
  wire  mem_0_65_W0_en;
  wire  mem_0_65_W0_mask;
  wire [6:0] mem_0_65_R0_addr;
  wire  mem_0_65_R0_clk;
  wire [7:0] mem_0_65_R0_data;
  wire  mem_0_65_R0_en;
  wire [6:0] mem_0_66_W0_addr;
  wire  mem_0_66_W0_clk;
  wire [7:0] mem_0_66_W0_data;
  wire  mem_0_66_W0_en;
  wire  mem_0_66_W0_mask;
  wire [6:0] mem_0_66_R0_addr;
  wire  mem_0_66_R0_clk;
  wire [7:0] mem_0_66_R0_data;
  wire  mem_0_66_R0_en;
  wire [6:0] mem_0_67_W0_addr;
  wire  mem_0_67_W0_clk;
  wire [7:0] mem_0_67_W0_data;
  wire  mem_0_67_W0_en;
  wire  mem_0_67_W0_mask;
  wire [6:0] mem_0_67_R0_addr;
  wire  mem_0_67_R0_clk;
  wire [7:0] mem_0_67_R0_data;
  wire  mem_0_67_R0_en;
  wire [6:0] mem_0_68_W0_addr;
  wire  mem_0_68_W0_clk;
  wire [7:0] mem_0_68_W0_data;
  wire  mem_0_68_W0_en;
  wire  mem_0_68_W0_mask;
  wire [6:0] mem_0_68_R0_addr;
  wire  mem_0_68_R0_clk;
  wire [7:0] mem_0_68_R0_data;
  wire  mem_0_68_R0_en;
  wire [6:0] mem_0_69_W0_addr;
  wire  mem_0_69_W0_clk;
  wire [7:0] mem_0_69_W0_data;
  wire  mem_0_69_W0_en;
  wire  mem_0_69_W0_mask;
  wire [6:0] mem_0_69_R0_addr;
  wire  mem_0_69_R0_clk;
  wire [7:0] mem_0_69_R0_data;
  wire  mem_0_69_R0_en;
  wire [6:0] mem_0_70_W0_addr;
  wire  mem_0_70_W0_clk;
  wire [7:0] mem_0_70_W0_data;
  wire  mem_0_70_W0_en;
  wire  mem_0_70_W0_mask;
  wire [6:0] mem_0_70_R0_addr;
  wire  mem_0_70_R0_clk;
  wire [7:0] mem_0_70_R0_data;
  wire  mem_0_70_R0_en;
  wire [6:0] mem_0_71_W0_addr;
  wire  mem_0_71_W0_clk;
  wire [7:0] mem_0_71_W0_data;
  wire  mem_0_71_W0_en;
  wire  mem_0_71_W0_mask;
  wire [6:0] mem_0_71_R0_addr;
  wire  mem_0_71_R0_clk;
  wire [7:0] mem_0_71_R0_data;
  wire  mem_0_71_R0_en;
  wire [6:0] mem_0_72_W0_addr;
  wire  mem_0_72_W0_clk;
  wire [7:0] mem_0_72_W0_data;
  wire  mem_0_72_W0_en;
  wire  mem_0_72_W0_mask;
  wire [6:0] mem_0_72_R0_addr;
  wire  mem_0_72_R0_clk;
  wire [7:0] mem_0_72_R0_data;
  wire  mem_0_72_R0_en;
  wire [6:0] mem_0_73_W0_addr;
  wire  mem_0_73_W0_clk;
  wire [7:0] mem_0_73_W0_data;
  wire  mem_0_73_W0_en;
  wire  mem_0_73_W0_mask;
  wire [6:0] mem_0_73_R0_addr;
  wire  mem_0_73_R0_clk;
  wire [7:0] mem_0_73_R0_data;
  wire  mem_0_73_R0_en;
  wire [6:0] mem_0_74_W0_addr;
  wire  mem_0_74_W0_clk;
  wire [7:0] mem_0_74_W0_data;
  wire  mem_0_74_W0_en;
  wire  mem_0_74_W0_mask;
  wire [6:0] mem_0_74_R0_addr;
  wire  mem_0_74_R0_clk;
  wire [7:0] mem_0_74_R0_data;
  wire  mem_0_74_R0_en;
  wire [6:0] mem_0_75_W0_addr;
  wire  mem_0_75_W0_clk;
  wire [7:0] mem_0_75_W0_data;
  wire  mem_0_75_W0_en;
  wire  mem_0_75_W0_mask;
  wire [6:0] mem_0_75_R0_addr;
  wire  mem_0_75_R0_clk;
  wire [7:0] mem_0_75_R0_data;
  wire  mem_0_75_R0_en;
  wire [6:0] mem_0_76_W0_addr;
  wire  mem_0_76_W0_clk;
  wire [7:0] mem_0_76_W0_data;
  wire  mem_0_76_W0_en;
  wire  mem_0_76_W0_mask;
  wire [6:0] mem_0_76_R0_addr;
  wire  mem_0_76_R0_clk;
  wire [7:0] mem_0_76_R0_data;
  wire  mem_0_76_R0_en;
  wire [6:0] mem_0_77_W0_addr;
  wire  mem_0_77_W0_clk;
  wire [7:0] mem_0_77_W0_data;
  wire  mem_0_77_W0_en;
  wire  mem_0_77_W0_mask;
  wire [6:0] mem_0_77_R0_addr;
  wire  mem_0_77_R0_clk;
  wire [7:0] mem_0_77_R0_data;
  wire  mem_0_77_R0_en;
  wire [6:0] mem_0_78_W0_addr;
  wire  mem_0_78_W0_clk;
  wire [7:0] mem_0_78_W0_data;
  wire  mem_0_78_W0_en;
  wire  mem_0_78_W0_mask;
  wire [6:0] mem_0_78_R0_addr;
  wire  mem_0_78_R0_clk;
  wire [7:0] mem_0_78_R0_data;
  wire  mem_0_78_R0_en;
  wire [6:0] mem_0_79_W0_addr;
  wire  mem_0_79_W0_clk;
  wire [7:0] mem_0_79_W0_data;
  wire  mem_0_79_W0_en;
  wire  mem_0_79_W0_mask;
  wire [6:0] mem_0_79_R0_addr;
  wire  mem_0_79_R0_clk;
  wire [7:0] mem_0_79_R0_data;
  wire  mem_0_79_R0_en;
  wire [6:0] mem_0_80_W0_addr;
  wire  mem_0_80_W0_clk;
  wire [7:0] mem_0_80_W0_data;
  wire  mem_0_80_W0_en;
  wire  mem_0_80_W0_mask;
  wire [6:0] mem_0_80_R0_addr;
  wire  mem_0_80_R0_clk;
  wire [7:0] mem_0_80_R0_data;
  wire  mem_0_80_R0_en;
  wire [6:0] mem_0_81_W0_addr;
  wire  mem_0_81_W0_clk;
  wire [7:0] mem_0_81_W0_data;
  wire  mem_0_81_W0_en;
  wire  mem_0_81_W0_mask;
  wire [6:0] mem_0_81_R0_addr;
  wire  mem_0_81_R0_clk;
  wire [7:0] mem_0_81_R0_data;
  wire  mem_0_81_R0_en;
  wire [6:0] mem_0_82_W0_addr;
  wire  mem_0_82_W0_clk;
  wire [7:0] mem_0_82_W0_data;
  wire  mem_0_82_W0_en;
  wire  mem_0_82_W0_mask;
  wire [6:0] mem_0_82_R0_addr;
  wire  mem_0_82_R0_clk;
  wire [7:0] mem_0_82_R0_data;
  wire  mem_0_82_R0_en;
  wire [6:0] mem_0_83_W0_addr;
  wire  mem_0_83_W0_clk;
  wire [7:0] mem_0_83_W0_data;
  wire  mem_0_83_W0_en;
  wire  mem_0_83_W0_mask;
  wire [6:0] mem_0_83_R0_addr;
  wire  mem_0_83_R0_clk;
  wire [7:0] mem_0_83_R0_data;
  wire  mem_0_83_R0_en;
  wire [6:0] mem_0_84_W0_addr;
  wire  mem_0_84_W0_clk;
  wire [7:0] mem_0_84_W0_data;
  wire  mem_0_84_W0_en;
  wire  mem_0_84_W0_mask;
  wire [6:0] mem_0_84_R0_addr;
  wire  mem_0_84_R0_clk;
  wire [7:0] mem_0_84_R0_data;
  wire  mem_0_84_R0_en;
  wire [6:0] mem_0_85_W0_addr;
  wire  mem_0_85_W0_clk;
  wire [7:0] mem_0_85_W0_data;
  wire  mem_0_85_W0_en;
  wire  mem_0_85_W0_mask;
  wire [6:0] mem_0_85_R0_addr;
  wire  mem_0_85_R0_clk;
  wire [7:0] mem_0_85_R0_data;
  wire  mem_0_85_R0_en;
  wire [6:0] mem_0_86_W0_addr;
  wire  mem_0_86_W0_clk;
  wire [7:0] mem_0_86_W0_data;
  wire  mem_0_86_W0_en;
  wire  mem_0_86_W0_mask;
  wire [6:0] mem_0_86_R0_addr;
  wire  mem_0_86_R0_clk;
  wire [7:0] mem_0_86_R0_data;
  wire  mem_0_86_R0_en;
  wire [6:0] mem_0_87_W0_addr;
  wire  mem_0_87_W0_clk;
  wire [7:0] mem_0_87_W0_data;
  wire  mem_0_87_W0_en;
  wire  mem_0_87_W0_mask;
  wire [6:0] mem_0_87_R0_addr;
  wire  mem_0_87_R0_clk;
  wire [7:0] mem_0_87_R0_data;
  wire  mem_0_87_R0_en;
  wire [6:0] mem_0_88_W0_addr;
  wire  mem_0_88_W0_clk;
  wire [7:0] mem_0_88_W0_data;
  wire  mem_0_88_W0_en;
  wire  mem_0_88_W0_mask;
  wire [6:0] mem_0_88_R0_addr;
  wire  mem_0_88_R0_clk;
  wire [7:0] mem_0_88_R0_data;
  wire  mem_0_88_R0_en;
  wire [6:0] mem_0_89_W0_addr;
  wire  mem_0_89_W0_clk;
  wire [7:0] mem_0_89_W0_data;
  wire  mem_0_89_W0_en;
  wire  mem_0_89_W0_mask;
  wire [6:0] mem_0_89_R0_addr;
  wire  mem_0_89_R0_clk;
  wire [7:0] mem_0_89_R0_data;
  wire  mem_0_89_R0_en;
  wire [6:0] mem_0_90_W0_addr;
  wire  mem_0_90_W0_clk;
  wire [7:0] mem_0_90_W0_data;
  wire  mem_0_90_W0_en;
  wire  mem_0_90_W0_mask;
  wire [6:0] mem_0_90_R0_addr;
  wire  mem_0_90_R0_clk;
  wire [7:0] mem_0_90_R0_data;
  wire  mem_0_90_R0_en;
  wire [6:0] mem_0_91_W0_addr;
  wire  mem_0_91_W0_clk;
  wire [7:0] mem_0_91_W0_data;
  wire  mem_0_91_W0_en;
  wire  mem_0_91_W0_mask;
  wire [6:0] mem_0_91_R0_addr;
  wire  mem_0_91_R0_clk;
  wire [7:0] mem_0_91_R0_data;
  wire  mem_0_91_R0_en;
  wire [6:0] mem_0_92_W0_addr;
  wire  mem_0_92_W0_clk;
  wire [7:0] mem_0_92_W0_data;
  wire  mem_0_92_W0_en;
  wire  mem_0_92_W0_mask;
  wire [6:0] mem_0_92_R0_addr;
  wire  mem_0_92_R0_clk;
  wire [7:0] mem_0_92_R0_data;
  wire  mem_0_92_R0_en;
  wire [6:0] mem_0_93_W0_addr;
  wire  mem_0_93_W0_clk;
  wire [7:0] mem_0_93_W0_data;
  wire  mem_0_93_W0_en;
  wire  mem_0_93_W0_mask;
  wire [6:0] mem_0_93_R0_addr;
  wire  mem_0_93_R0_clk;
  wire [7:0] mem_0_93_R0_data;
  wire  mem_0_93_R0_en;
  wire [6:0] mem_0_94_W0_addr;
  wire  mem_0_94_W0_clk;
  wire [7:0] mem_0_94_W0_data;
  wire  mem_0_94_W0_en;
  wire  mem_0_94_W0_mask;
  wire [6:0] mem_0_94_R0_addr;
  wire  mem_0_94_R0_clk;
  wire [7:0] mem_0_94_R0_data;
  wire  mem_0_94_R0_en;
  wire [6:0] mem_0_95_W0_addr;
  wire  mem_0_95_W0_clk;
  wire [7:0] mem_0_95_W0_data;
  wire  mem_0_95_W0_en;
  wire  mem_0_95_W0_mask;
  wire [6:0] mem_0_95_R0_addr;
  wire  mem_0_95_R0_clk;
  wire [7:0] mem_0_95_R0_data;
  wire  mem_0_95_R0_en;
  wire [6:0] mem_0_96_W0_addr;
  wire  mem_0_96_W0_clk;
  wire [7:0] mem_0_96_W0_data;
  wire  mem_0_96_W0_en;
  wire  mem_0_96_W0_mask;
  wire [6:0] mem_0_96_R0_addr;
  wire  mem_0_96_R0_clk;
  wire [7:0] mem_0_96_R0_data;
  wire  mem_0_96_R0_en;
  wire [6:0] mem_0_97_W0_addr;
  wire  mem_0_97_W0_clk;
  wire [7:0] mem_0_97_W0_data;
  wire  mem_0_97_W0_en;
  wire  mem_0_97_W0_mask;
  wire [6:0] mem_0_97_R0_addr;
  wire  mem_0_97_R0_clk;
  wire [7:0] mem_0_97_R0_data;
  wire  mem_0_97_R0_en;
  wire [6:0] mem_0_98_W0_addr;
  wire  mem_0_98_W0_clk;
  wire [7:0] mem_0_98_W0_data;
  wire  mem_0_98_W0_en;
  wire  mem_0_98_W0_mask;
  wire [6:0] mem_0_98_R0_addr;
  wire  mem_0_98_R0_clk;
  wire [7:0] mem_0_98_R0_data;
  wire  mem_0_98_R0_en;
  wire [6:0] mem_0_99_W0_addr;
  wire  mem_0_99_W0_clk;
  wire [7:0] mem_0_99_W0_data;
  wire  mem_0_99_W0_en;
  wire  mem_0_99_W0_mask;
  wire [6:0] mem_0_99_R0_addr;
  wire  mem_0_99_R0_clk;
  wire [7:0] mem_0_99_R0_data;
  wire  mem_0_99_R0_en;
  wire [6:0] mem_0_100_W0_addr;
  wire  mem_0_100_W0_clk;
  wire [7:0] mem_0_100_W0_data;
  wire  mem_0_100_W0_en;
  wire  mem_0_100_W0_mask;
  wire [6:0] mem_0_100_R0_addr;
  wire  mem_0_100_R0_clk;
  wire [7:0] mem_0_100_R0_data;
  wire  mem_0_100_R0_en;
  wire [6:0] mem_0_101_W0_addr;
  wire  mem_0_101_W0_clk;
  wire [7:0] mem_0_101_W0_data;
  wire  mem_0_101_W0_en;
  wire  mem_0_101_W0_mask;
  wire [6:0] mem_0_101_R0_addr;
  wire  mem_0_101_R0_clk;
  wire [7:0] mem_0_101_R0_data;
  wire  mem_0_101_R0_en;
  wire [6:0] mem_0_102_W0_addr;
  wire  mem_0_102_W0_clk;
  wire [7:0] mem_0_102_W0_data;
  wire  mem_0_102_W0_en;
  wire  mem_0_102_W0_mask;
  wire [6:0] mem_0_102_R0_addr;
  wire  mem_0_102_R0_clk;
  wire [7:0] mem_0_102_R0_data;
  wire  mem_0_102_R0_en;
  wire [6:0] mem_0_103_W0_addr;
  wire  mem_0_103_W0_clk;
  wire [7:0] mem_0_103_W0_data;
  wire  mem_0_103_W0_en;
  wire  mem_0_103_W0_mask;
  wire [6:0] mem_0_103_R0_addr;
  wire  mem_0_103_R0_clk;
  wire [7:0] mem_0_103_R0_data;
  wire  mem_0_103_R0_en;
  wire [6:0] mem_0_104_W0_addr;
  wire  mem_0_104_W0_clk;
  wire [7:0] mem_0_104_W0_data;
  wire  mem_0_104_W0_en;
  wire  mem_0_104_W0_mask;
  wire [6:0] mem_0_104_R0_addr;
  wire  mem_0_104_R0_clk;
  wire [7:0] mem_0_104_R0_data;
  wire  mem_0_104_R0_en;
  wire [6:0] mem_0_105_W0_addr;
  wire  mem_0_105_W0_clk;
  wire [7:0] mem_0_105_W0_data;
  wire  mem_0_105_W0_en;
  wire  mem_0_105_W0_mask;
  wire [6:0] mem_0_105_R0_addr;
  wire  mem_0_105_R0_clk;
  wire [7:0] mem_0_105_R0_data;
  wire  mem_0_105_R0_en;
  wire [6:0] mem_0_106_W0_addr;
  wire  mem_0_106_W0_clk;
  wire [7:0] mem_0_106_W0_data;
  wire  mem_0_106_W0_en;
  wire  mem_0_106_W0_mask;
  wire [6:0] mem_0_106_R0_addr;
  wire  mem_0_106_R0_clk;
  wire [7:0] mem_0_106_R0_data;
  wire  mem_0_106_R0_en;
  wire [6:0] mem_0_107_W0_addr;
  wire  mem_0_107_W0_clk;
  wire [7:0] mem_0_107_W0_data;
  wire  mem_0_107_W0_en;
  wire  mem_0_107_W0_mask;
  wire [6:0] mem_0_107_R0_addr;
  wire  mem_0_107_R0_clk;
  wire [7:0] mem_0_107_R0_data;
  wire  mem_0_107_R0_en;
  wire [6:0] mem_0_108_W0_addr;
  wire  mem_0_108_W0_clk;
  wire [7:0] mem_0_108_W0_data;
  wire  mem_0_108_W0_en;
  wire  mem_0_108_W0_mask;
  wire [6:0] mem_0_108_R0_addr;
  wire  mem_0_108_R0_clk;
  wire [7:0] mem_0_108_R0_data;
  wire  mem_0_108_R0_en;
  wire [6:0] mem_0_109_W0_addr;
  wire  mem_0_109_W0_clk;
  wire [7:0] mem_0_109_W0_data;
  wire  mem_0_109_W0_en;
  wire  mem_0_109_W0_mask;
  wire [6:0] mem_0_109_R0_addr;
  wire  mem_0_109_R0_clk;
  wire [7:0] mem_0_109_R0_data;
  wire  mem_0_109_R0_en;
  wire [6:0] mem_0_110_W0_addr;
  wire  mem_0_110_W0_clk;
  wire [7:0] mem_0_110_W0_data;
  wire  mem_0_110_W0_en;
  wire  mem_0_110_W0_mask;
  wire [6:0] mem_0_110_R0_addr;
  wire  mem_0_110_R0_clk;
  wire [7:0] mem_0_110_R0_data;
  wire  mem_0_110_R0_en;
  wire [6:0] mem_0_111_W0_addr;
  wire  mem_0_111_W0_clk;
  wire [7:0] mem_0_111_W0_data;
  wire  mem_0_111_W0_en;
  wire  mem_0_111_W0_mask;
  wire [6:0] mem_0_111_R0_addr;
  wire  mem_0_111_R0_clk;
  wire [7:0] mem_0_111_R0_data;
  wire  mem_0_111_R0_en;
  wire [6:0] mem_0_112_W0_addr;
  wire  mem_0_112_W0_clk;
  wire [7:0] mem_0_112_W0_data;
  wire  mem_0_112_W0_en;
  wire  mem_0_112_W0_mask;
  wire [6:0] mem_0_112_R0_addr;
  wire  mem_0_112_R0_clk;
  wire [7:0] mem_0_112_R0_data;
  wire  mem_0_112_R0_en;
  wire [6:0] mem_0_113_W0_addr;
  wire  mem_0_113_W0_clk;
  wire [7:0] mem_0_113_W0_data;
  wire  mem_0_113_W0_en;
  wire  mem_0_113_W0_mask;
  wire [6:0] mem_0_113_R0_addr;
  wire  mem_0_113_R0_clk;
  wire [7:0] mem_0_113_R0_data;
  wire  mem_0_113_R0_en;
  wire [6:0] mem_0_114_W0_addr;
  wire  mem_0_114_W0_clk;
  wire [7:0] mem_0_114_W0_data;
  wire  mem_0_114_W0_en;
  wire  mem_0_114_W0_mask;
  wire [6:0] mem_0_114_R0_addr;
  wire  mem_0_114_R0_clk;
  wire [7:0] mem_0_114_R0_data;
  wire  mem_0_114_R0_en;
  wire [6:0] mem_0_115_W0_addr;
  wire  mem_0_115_W0_clk;
  wire [7:0] mem_0_115_W0_data;
  wire  mem_0_115_W0_en;
  wire  mem_0_115_W0_mask;
  wire [6:0] mem_0_115_R0_addr;
  wire  mem_0_115_R0_clk;
  wire [7:0] mem_0_115_R0_data;
  wire  mem_0_115_R0_en;
  wire [6:0] mem_0_116_W0_addr;
  wire  mem_0_116_W0_clk;
  wire [7:0] mem_0_116_W0_data;
  wire  mem_0_116_W0_en;
  wire  mem_0_116_W0_mask;
  wire [6:0] mem_0_116_R0_addr;
  wire  mem_0_116_R0_clk;
  wire [7:0] mem_0_116_R0_data;
  wire  mem_0_116_R0_en;
  wire [6:0] mem_0_117_W0_addr;
  wire  mem_0_117_W0_clk;
  wire [7:0] mem_0_117_W0_data;
  wire  mem_0_117_W0_en;
  wire  mem_0_117_W0_mask;
  wire [6:0] mem_0_117_R0_addr;
  wire  mem_0_117_R0_clk;
  wire [7:0] mem_0_117_R0_data;
  wire  mem_0_117_R0_en;
  wire [6:0] mem_0_118_W0_addr;
  wire  mem_0_118_W0_clk;
  wire [7:0] mem_0_118_W0_data;
  wire  mem_0_118_W0_en;
  wire  mem_0_118_W0_mask;
  wire [6:0] mem_0_118_R0_addr;
  wire  mem_0_118_R0_clk;
  wire [7:0] mem_0_118_R0_data;
  wire  mem_0_118_R0_en;
  wire [6:0] mem_0_119_W0_addr;
  wire  mem_0_119_W0_clk;
  wire [7:0] mem_0_119_W0_data;
  wire  mem_0_119_W0_en;
  wire  mem_0_119_W0_mask;
  wire [6:0] mem_0_119_R0_addr;
  wire  mem_0_119_R0_clk;
  wire [7:0] mem_0_119_R0_data;
  wire  mem_0_119_R0_en;
  wire [6:0] mem_0_120_W0_addr;
  wire  mem_0_120_W0_clk;
  wire [7:0] mem_0_120_W0_data;
  wire  mem_0_120_W0_en;
  wire  mem_0_120_W0_mask;
  wire [6:0] mem_0_120_R0_addr;
  wire  mem_0_120_R0_clk;
  wire [7:0] mem_0_120_R0_data;
  wire  mem_0_120_R0_en;
  wire [6:0] mem_0_121_W0_addr;
  wire  mem_0_121_W0_clk;
  wire [7:0] mem_0_121_W0_data;
  wire  mem_0_121_W0_en;
  wire  mem_0_121_W0_mask;
  wire [6:0] mem_0_121_R0_addr;
  wire  mem_0_121_R0_clk;
  wire [7:0] mem_0_121_R0_data;
  wire  mem_0_121_R0_en;
  wire [6:0] mem_0_122_W0_addr;
  wire  mem_0_122_W0_clk;
  wire [7:0] mem_0_122_W0_data;
  wire  mem_0_122_W0_en;
  wire  mem_0_122_W0_mask;
  wire [6:0] mem_0_122_R0_addr;
  wire  mem_0_122_R0_clk;
  wire [7:0] mem_0_122_R0_data;
  wire  mem_0_122_R0_en;
  wire [6:0] mem_0_123_W0_addr;
  wire  mem_0_123_W0_clk;
  wire [7:0] mem_0_123_W0_data;
  wire  mem_0_123_W0_en;
  wire  mem_0_123_W0_mask;
  wire [6:0] mem_0_123_R0_addr;
  wire  mem_0_123_R0_clk;
  wire [7:0] mem_0_123_R0_data;
  wire  mem_0_123_R0_en;
  wire [6:0] mem_0_124_W0_addr;
  wire  mem_0_124_W0_clk;
  wire [7:0] mem_0_124_W0_data;
  wire  mem_0_124_W0_en;
  wire  mem_0_124_W0_mask;
  wire [6:0] mem_0_124_R0_addr;
  wire  mem_0_124_R0_clk;
  wire [7:0] mem_0_124_R0_data;
  wire  mem_0_124_R0_en;
  wire [6:0] mem_0_125_W0_addr;
  wire  mem_0_125_W0_clk;
  wire [7:0] mem_0_125_W0_data;
  wire  mem_0_125_W0_en;
  wire  mem_0_125_W0_mask;
  wire [6:0] mem_0_125_R0_addr;
  wire  mem_0_125_R0_clk;
  wire [7:0] mem_0_125_R0_data;
  wire  mem_0_125_R0_en;
  wire [6:0] mem_0_126_W0_addr;
  wire  mem_0_126_W0_clk;
  wire [7:0] mem_0_126_W0_data;
  wire  mem_0_126_W0_en;
  wire  mem_0_126_W0_mask;
  wire [6:0] mem_0_126_R0_addr;
  wire  mem_0_126_R0_clk;
  wire [7:0] mem_0_126_R0_data;
  wire  mem_0_126_R0_en;
  wire [6:0] mem_0_127_W0_addr;
  wire  mem_0_127_W0_clk;
  wire [7:0] mem_0_127_W0_data;
  wire  mem_0_127_W0_en;
  wire  mem_0_127_W0_mask;
  wire [6:0] mem_0_127_R0_addr;
  wire  mem_0_127_R0_clk;
  wire [7:0] mem_0_127_R0_data;
  wire  mem_0_127_R0_en;
  wire [6:0] mem_0_128_W0_addr;
  wire  mem_0_128_W0_clk;
  wire [7:0] mem_0_128_W0_data;
  wire  mem_0_128_W0_en;
  wire  mem_0_128_W0_mask;
  wire [6:0] mem_0_128_R0_addr;
  wire  mem_0_128_R0_clk;
  wire [7:0] mem_0_128_R0_data;
  wire  mem_0_128_R0_en;
  wire [6:0] mem_0_129_W0_addr;
  wire  mem_0_129_W0_clk;
  wire [7:0] mem_0_129_W0_data;
  wire  mem_0_129_W0_en;
  wire  mem_0_129_W0_mask;
  wire [6:0] mem_0_129_R0_addr;
  wire  mem_0_129_R0_clk;
  wire [7:0] mem_0_129_R0_data;
  wire  mem_0_129_R0_en;
  wire [6:0] mem_0_130_W0_addr;
  wire  mem_0_130_W0_clk;
  wire [7:0] mem_0_130_W0_data;
  wire  mem_0_130_W0_en;
  wire  mem_0_130_W0_mask;
  wire [6:0] mem_0_130_R0_addr;
  wire  mem_0_130_R0_clk;
  wire [7:0] mem_0_130_R0_data;
  wire  mem_0_130_R0_en;
  wire [6:0] mem_0_131_W0_addr;
  wire  mem_0_131_W0_clk;
  wire [7:0] mem_0_131_W0_data;
  wire  mem_0_131_W0_en;
  wire  mem_0_131_W0_mask;
  wire [6:0] mem_0_131_R0_addr;
  wire  mem_0_131_R0_clk;
  wire [7:0] mem_0_131_R0_data;
  wire  mem_0_131_R0_en;
  wire [6:0] mem_0_132_W0_addr;
  wire  mem_0_132_W0_clk;
  wire [7:0] mem_0_132_W0_data;
  wire  mem_0_132_W0_en;
  wire  mem_0_132_W0_mask;
  wire [6:0] mem_0_132_R0_addr;
  wire  mem_0_132_R0_clk;
  wire [7:0] mem_0_132_R0_data;
  wire  mem_0_132_R0_en;
  wire [6:0] mem_0_133_W0_addr;
  wire  mem_0_133_W0_clk;
  wire [7:0] mem_0_133_W0_data;
  wire  mem_0_133_W0_en;
  wire  mem_0_133_W0_mask;
  wire [6:0] mem_0_133_R0_addr;
  wire  mem_0_133_R0_clk;
  wire [7:0] mem_0_133_R0_data;
  wire  mem_0_133_R0_en;
  wire [6:0] mem_0_134_W0_addr;
  wire  mem_0_134_W0_clk;
  wire [7:0] mem_0_134_W0_data;
  wire  mem_0_134_W0_en;
  wire  mem_0_134_W0_mask;
  wire [6:0] mem_0_134_R0_addr;
  wire  mem_0_134_R0_clk;
  wire [7:0] mem_0_134_R0_data;
  wire  mem_0_134_R0_en;
  wire [6:0] mem_0_135_W0_addr;
  wire  mem_0_135_W0_clk;
  wire [7:0] mem_0_135_W0_data;
  wire  mem_0_135_W0_en;
  wire  mem_0_135_W0_mask;
  wire [6:0] mem_0_135_R0_addr;
  wire  mem_0_135_R0_clk;
  wire [7:0] mem_0_135_R0_data;
  wire  mem_0_135_R0_en;
  wire [6:0] mem_0_136_W0_addr;
  wire  mem_0_136_W0_clk;
  wire [7:0] mem_0_136_W0_data;
  wire  mem_0_136_W0_en;
  wire  mem_0_136_W0_mask;
  wire [6:0] mem_0_136_R0_addr;
  wire  mem_0_136_R0_clk;
  wire [7:0] mem_0_136_R0_data;
  wire  mem_0_136_R0_en;
  wire [6:0] mem_0_137_W0_addr;
  wire  mem_0_137_W0_clk;
  wire [7:0] mem_0_137_W0_data;
  wire  mem_0_137_W0_en;
  wire  mem_0_137_W0_mask;
  wire [6:0] mem_0_137_R0_addr;
  wire  mem_0_137_R0_clk;
  wire [7:0] mem_0_137_R0_data;
  wire  mem_0_137_R0_en;
  wire [6:0] mem_0_138_W0_addr;
  wire  mem_0_138_W0_clk;
  wire [7:0] mem_0_138_W0_data;
  wire  mem_0_138_W0_en;
  wire  mem_0_138_W0_mask;
  wire [6:0] mem_0_138_R0_addr;
  wire  mem_0_138_R0_clk;
  wire [7:0] mem_0_138_R0_data;
  wire  mem_0_138_R0_en;
  wire [6:0] mem_0_139_W0_addr;
  wire  mem_0_139_W0_clk;
  wire [7:0] mem_0_139_W0_data;
  wire  mem_0_139_W0_en;
  wire  mem_0_139_W0_mask;
  wire [6:0] mem_0_139_R0_addr;
  wire  mem_0_139_R0_clk;
  wire [7:0] mem_0_139_R0_data;
  wire  mem_0_139_R0_en;
  wire [6:0] mem_0_140_W0_addr;
  wire  mem_0_140_W0_clk;
  wire [7:0] mem_0_140_W0_data;
  wire  mem_0_140_W0_en;
  wire  mem_0_140_W0_mask;
  wire [6:0] mem_0_140_R0_addr;
  wire  mem_0_140_R0_clk;
  wire [7:0] mem_0_140_R0_data;
  wire  mem_0_140_R0_en;
  wire [6:0] mem_0_141_W0_addr;
  wire  mem_0_141_W0_clk;
  wire [7:0] mem_0_141_W0_data;
  wire  mem_0_141_W0_en;
  wire  mem_0_141_W0_mask;
  wire [6:0] mem_0_141_R0_addr;
  wire  mem_0_141_R0_clk;
  wire [7:0] mem_0_141_R0_data;
  wire  mem_0_141_R0_en;
  wire [6:0] mem_0_142_W0_addr;
  wire  mem_0_142_W0_clk;
  wire [7:0] mem_0_142_W0_data;
  wire  mem_0_142_W0_en;
  wire  mem_0_142_W0_mask;
  wire [6:0] mem_0_142_R0_addr;
  wire  mem_0_142_R0_clk;
  wire [7:0] mem_0_142_R0_data;
  wire  mem_0_142_R0_en;
  wire [6:0] mem_0_143_W0_addr;
  wire  mem_0_143_W0_clk;
  wire [7:0] mem_0_143_W0_data;
  wire  mem_0_143_W0_en;
  wire  mem_0_143_W0_mask;
  wire [6:0] mem_0_143_R0_addr;
  wire  mem_0_143_R0_clk;
  wire [7:0] mem_0_143_R0_data;
  wire  mem_0_143_R0_en;
  wire [6:0] mem_0_144_W0_addr;
  wire  mem_0_144_W0_clk;
  wire [7:0] mem_0_144_W0_data;
  wire  mem_0_144_W0_en;
  wire  mem_0_144_W0_mask;
  wire [6:0] mem_0_144_R0_addr;
  wire  mem_0_144_R0_clk;
  wire [7:0] mem_0_144_R0_data;
  wire  mem_0_144_R0_en;
  wire [6:0] mem_0_145_W0_addr;
  wire  mem_0_145_W0_clk;
  wire [7:0] mem_0_145_W0_data;
  wire  mem_0_145_W0_en;
  wire  mem_0_145_W0_mask;
  wire [6:0] mem_0_145_R0_addr;
  wire  mem_0_145_R0_clk;
  wire [7:0] mem_0_145_R0_data;
  wire  mem_0_145_R0_en;
  wire [6:0] mem_0_146_W0_addr;
  wire  mem_0_146_W0_clk;
  wire [7:0] mem_0_146_W0_data;
  wire  mem_0_146_W0_en;
  wire  mem_0_146_W0_mask;
  wire [6:0] mem_0_146_R0_addr;
  wire  mem_0_146_R0_clk;
  wire [7:0] mem_0_146_R0_data;
  wire  mem_0_146_R0_en;
  wire [6:0] mem_0_147_W0_addr;
  wire  mem_0_147_W0_clk;
  wire [7:0] mem_0_147_W0_data;
  wire  mem_0_147_W0_en;
  wire  mem_0_147_W0_mask;
  wire [6:0] mem_0_147_R0_addr;
  wire  mem_0_147_R0_clk;
  wire [7:0] mem_0_147_R0_data;
  wire  mem_0_147_R0_en;
  wire [6:0] mem_0_148_W0_addr;
  wire  mem_0_148_W0_clk;
  wire [7:0] mem_0_148_W0_data;
  wire  mem_0_148_W0_en;
  wire  mem_0_148_W0_mask;
  wire [6:0] mem_0_148_R0_addr;
  wire  mem_0_148_R0_clk;
  wire [7:0] mem_0_148_R0_data;
  wire  mem_0_148_R0_en;
  wire [6:0] mem_0_149_W0_addr;
  wire  mem_0_149_W0_clk;
  wire [7:0] mem_0_149_W0_data;
  wire  mem_0_149_W0_en;
  wire  mem_0_149_W0_mask;
  wire [6:0] mem_0_149_R0_addr;
  wire  mem_0_149_R0_clk;
  wire [7:0] mem_0_149_R0_data;
  wire  mem_0_149_R0_en;
  wire [6:0] mem_0_150_W0_addr;
  wire  mem_0_150_W0_clk;
  wire [7:0] mem_0_150_W0_data;
  wire  mem_0_150_W0_en;
  wire  mem_0_150_W0_mask;
  wire [6:0] mem_0_150_R0_addr;
  wire  mem_0_150_R0_clk;
  wire [7:0] mem_0_150_R0_data;
  wire  mem_0_150_R0_en;
  wire [6:0] mem_0_151_W0_addr;
  wire  mem_0_151_W0_clk;
  wire [7:0] mem_0_151_W0_data;
  wire  mem_0_151_W0_en;
  wire  mem_0_151_W0_mask;
  wire [6:0] mem_0_151_R0_addr;
  wire  mem_0_151_R0_clk;
  wire [7:0] mem_0_151_R0_data;
  wire  mem_0_151_R0_en;
  wire [6:0] mem_0_152_W0_addr;
  wire  mem_0_152_W0_clk;
  wire [7:0] mem_0_152_W0_data;
  wire  mem_0_152_W0_en;
  wire  mem_0_152_W0_mask;
  wire [6:0] mem_0_152_R0_addr;
  wire  mem_0_152_R0_clk;
  wire [7:0] mem_0_152_R0_data;
  wire  mem_0_152_R0_en;
  wire [6:0] mem_0_153_W0_addr;
  wire  mem_0_153_W0_clk;
  wire [7:0] mem_0_153_W0_data;
  wire  mem_0_153_W0_en;
  wire  mem_0_153_W0_mask;
  wire [6:0] mem_0_153_R0_addr;
  wire  mem_0_153_R0_clk;
  wire [7:0] mem_0_153_R0_data;
  wire  mem_0_153_R0_en;
  wire [6:0] mem_0_154_W0_addr;
  wire  mem_0_154_W0_clk;
  wire [7:0] mem_0_154_W0_data;
  wire  mem_0_154_W0_en;
  wire  mem_0_154_W0_mask;
  wire [6:0] mem_0_154_R0_addr;
  wire  mem_0_154_R0_clk;
  wire [7:0] mem_0_154_R0_data;
  wire  mem_0_154_R0_en;
  wire [6:0] mem_0_155_W0_addr;
  wire  mem_0_155_W0_clk;
  wire [7:0] mem_0_155_W0_data;
  wire  mem_0_155_W0_en;
  wire  mem_0_155_W0_mask;
  wire [6:0] mem_0_155_R0_addr;
  wire  mem_0_155_R0_clk;
  wire [7:0] mem_0_155_R0_data;
  wire  mem_0_155_R0_en;
  wire [6:0] mem_0_156_W0_addr;
  wire  mem_0_156_W0_clk;
  wire [7:0] mem_0_156_W0_data;
  wire  mem_0_156_W0_en;
  wire  mem_0_156_W0_mask;
  wire [6:0] mem_0_156_R0_addr;
  wire  mem_0_156_R0_clk;
  wire [7:0] mem_0_156_R0_data;
  wire  mem_0_156_R0_en;
  wire [6:0] mem_0_157_W0_addr;
  wire  mem_0_157_W0_clk;
  wire [7:0] mem_0_157_W0_data;
  wire  mem_0_157_W0_en;
  wire  mem_0_157_W0_mask;
  wire [6:0] mem_0_157_R0_addr;
  wire  mem_0_157_R0_clk;
  wire [7:0] mem_0_157_R0_data;
  wire  mem_0_157_R0_en;
  wire [6:0] mem_0_158_W0_addr;
  wire  mem_0_158_W0_clk;
  wire [7:0] mem_0_158_W0_data;
  wire  mem_0_158_W0_en;
  wire  mem_0_158_W0_mask;
  wire [6:0] mem_0_158_R0_addr;
  wire  mem_0_158_R0_clk;
  wire [7:0] mem_0_158_R0_data;
  wire  mem_0_158_R0_en;
  wire [6:0] mem_0_159_W0_addr;
  wire  mem_0_159_W0_clk;
  wire [7:0] mem_0_159_W0_data;
  wire  mem_0_159_W0_en;
  wire  mem_0_159_W0_mask;
  wire [6:0] mem_0_159_R0_addr;
  wire  mem_0_159_R0_clk;
  wire [7:0] mem_0_159_R0_data;
  wire  mem_0_159_R0_en;
  wire [6:0] mem_0_160_W0_addr;
  wire  mem_0_160_W0_clk;
  wire [7:0] mem_0_160_W0_data;
  wire  mem_0_160_W0_en;
  wire  mem_0_160_W0_mask;
  wire [6:0] mem_0_160_R0_addr;
  wire  mem_0_160_R0_clk;
  wire [7:0] mem_0_160_R0_data;
  wire  mem_0_160_R0_en;
  wire [6:0] mem_0_161_W0_addr;
  wire  mem_0_161_W0_clk;
  wire [7:0] mem_0_161_W0_data;
  wire  mem_0_161_W0_en;
  wire  mem_0_161_W0_mask;
  wire [6:0] mem_0_161_R0_addr;
  wire  mem_0_161_R0_clk;
  wire [7:0] mem_0_161_R0_data;
  wire  mem_0_161_R0_en;
  wire [6:0] mem_0_162_W0_addr;
  wire  mem_0_162_W0_clk;
  wire [7:0] mem_0_162_W0_data;
  wire  mem_0_162_W0_en;
  wire  mem_0_162_W0_mask;
  wire [6:0] mem_0_162_R0_addr;
  wire  mem_0_162_R0_clk;
  wire [7:0] mem_0_162_R0_data;
  wire  mem_0_162_R0_en;
  wire [6:0] mem_0_163_W0_addr;
  wire  mem_0_163_W0_clk;
  wire [7:0] mem_0_163_W0_data;
  wire  mem_0_163_W0_en;
  wire  mem_0_163_W0_mask;
  wire [6:0] mem_0_163_R0_addr;
  wire  mem_0_163_R0_clk;
  wire [7:0] mem_0_163_R0_data;
  wire  mem_0_163_R0_en;
  wire [6:0] mem_0_164_W0_addr;
  wire  mem_0_164_W0_clk;
  wire [7:0] mem_0_164_W0_data;
  wire  mem_0_164_W0_en;
  wire  mem_0_164_W0_mask;
  wire [6:0] mem_0_164_R0_addr;
  wire  mem_0_164_R0_clk;
  wire [7:0] mem_0_164_R0_data;
  wire  mem_0_164_R0_en;
  wire [6:0] mem_0_165_W0_addr;
  wire  mem_0_165_W0_clk;
  wire [7:0] mem_0_165_W0_data;
  wire  mem_0_165_W0_en;
  wire  mem_0_165_W0_mask;
  wire [6:0] mem_0_165_R0_addr;
  wire  mem_0_165_R0_clk;
  wire [7:0] mem_0_165_R0_data;
  wire  mem_0_165_R0_en;
  wire [6:0] mem_0_166_W0_addr;
  wire  mem_0_166_W0_clk;
  wire [7:0] mem_0_166_W0_data;
  wire  mem_0_166_W0_en;
  wire  mem_0_166_W0_mask;
  wire [6:0] mem_0_166_R0_addr;
  wire  mem_0_166_R0_clk;
  wire [7:0] mem_0_166_R0_data;
  wire  mem_0_166_R0_en;
  wire [6:0] mem_0_167_W0_addr;
  wire  mem_0_167_W0_clk;
  wire [7:0] mem_0_167_W0_data;
  wire  mem_0_167_W0_en;
  wire  mem_0_167_W0_mask;
  wire [6:0] mem_0_167_R0_addr;
  wire  mem_0_167_R0_clk;
  wire [7:0] mem_0_167_R0_data;
  wire  mem_0_167_R0_en;
  wire [6:0] mem_0_168_W0_addr;
  wire  mem_0_168_W0_clk;
  wire [7:0] mem_0_168_W0_data;
  wire  mem_0_168_W0_en;
  wire  mem_0_168_W0_mask;
  wire [6:0] mem_0_168_R0_addr;
  wire  mem_0_168_R0_clk;
  wire [7:0] mem_0_168_R0_data;
  wire  mem_0_168_R0_en;
  wire [6:0] mem_0_169_W0_addr;
  wire  mem_0_169_W0_clk;
  wire [7:0] mem_0_169_W0_data;
  wire  mem_0_169_W0_en;
  wire  mem_0_169_W0_mask;
  wire [6:0] mem_0_169_R0_addr;
  wire  mem_0_169_R0_clk;
  wire [7:0] mem_0_169_R0_data;
  wire  mem_0_169_R0_en;
  wire [6:0] mem_0_170_W0_addr;
  wire  mem_0_170_W0_clk;
  wire [7:0] mem_0_170_W0_data;
  wire  mem_0_170_W0_en;
  wire  mem_0_170_W0_mask;
  wire [6:0] mem_0_170_R0_addr;
  wire  mem_0_170_R0_clk;
  wire [7:0] mem_0_170_R0_data;
  wire  mem_0_170_R0_en;
  wire [6:0] mem_0_171_W0_addr;
  wire  mem_0_171_W0_clk;
  wire [7:0] mem_0_171_W0_data;
  wire  mem_0_171_W0_en;
  wire  mem_0_171_W0_mask;
  wire [6:0] mem_0_171_R0_addr;
  wire  mem_0_171_R0_clk;
  wire [7:0] mem_0_171_R0_data;
  wire  mem_0_171_R0_en;
  wire [6:0] mem_0_172_W0_addr;
  wire  mem_0_172_W0_clk;
  wire [7:0] mem_0_172_W0_data;
  wire  mem_0_172_W0_en;
  wire  mem_0_172_W0_mask;
  wire [6:0] mem_0_172_R0_addr;
  wire  mem_0_172_R0_clk;
  wire [7:0] mem_0_172_R0_data;
  wire  mem_0_172_R0_en;
  wire [6:0] mem_0_173_W0_addr;
  wire  mem_0_173_W0_clk;
  wire [7:0] mem_0_173_W0_data;
  wire  mem_0_173_W0_en;
  wire  mem_0_173_W0_mask;
  wire [6:0] mem_0_173_R0_addr;
  wire  mem_0_173_R0_clk;
  wire [7:0] mem_0_173_R0_data;
  wire  mem_0_173_R0_en;
  wire [6:0] mem_0_174_W0_addr;
  wire  mem_0_174_W0_clk;
  wire [7:0] mem_0_174_W0_data;
  wire  mem_0_174_W0_en;
  wire  mem_0_174_W0_mask;
  wire [6:0] mem_0_174_R0_addr;
  wire  mem_0_174_R0_clk;
  wire [7:0] mem_0_174_R0_data;
  wire  mem_0_174_R0_en;
  wire [6:0] mem_0_175_W0_addr;
  wire  mem_0_175_W0_clk;
  wire [7:0] mem_0_175_W0_data;
  wire  mem_0_175_W0_en;
  wire  mem_0_175_W0_mask;
  wire [6:0] mem_0_175_R0_addr;
  wire  mem_0_175_R0_clk;
  wire [7:0] mem_0_175_R0_data;
  wire  mem_0_175_R0_en;
  wire [6:0] mem_0_176_W0_addr;
  wire  mem_0_176_W0_clk;
  wire [7:0] mem_0_176_W0_data;
  wire  mem_0_176_W0_en;
  wire  mem_0_176_W0_mask;
  wire [6:0] mem_0_176_R0_addr;
  wire  mem_0_176_R0_clk;
  wire [7:0] mem_0_176_R0_data;
  wire  mem_0_176_R0_en;
  wire [6:0] mem_0_177_W0_addr;
  wire  mem_0_177_W0_clk;
  wire [7:0] mem_0_177_W0_data;
  wire  mem_0_177_W0_en;
  wire  mem_0_177_W0_mask;
  wire [6:0] mem_0_177_R0_addr;
  wire  mem_0_177_R0_clk;
  wire [7:0] mem_0_177_R0_data;
  wire  mem_0_177_R0_en;
  wire [6:0] mem_0_178_W0_addr;
  wire  mem_0_178_W0_clk;
  wire [7:0] mem_0_178_W0_data;
  wire  mem_0_178_W0_en;
  wire  mem_0_178_W0_mask;
  wire [6:0] mem_0_178_R0_addr;
  wire  mem_0_178_R0_clk;
  wire [7:0] mem_0_178_R0_data;
  wire  mem_0_178_R0_en;
  wire [6:0] mem_0_179_W0_addr;
  wire  mem_0_179_W0_clk;
  wire [7:0] mem_0_179_W0_data;
  wire  mem_0_179_W0_en;
  wire  mem_0_179_W0_mask;
  wire [6:0] mem_0_179_R0_addr;
  wire  mem_0_179_R0_clk;
  wire [7:0] mem_0_179_R0_data;
  wire  mem_0_179_R0_en;
  wire [6:0] mem_0_180_W0_addr;
  wire  mem_0_180_W0_clk;
  wire [7:0] mem_0_180_W0_data;
  wire  mem_0_180_W0_en;
  wire  mem_0_180_W0_mask;
  wire [6:0] mem_0_180_R0_addr;
  wire  mem_0_180_R0_clk;
  wire [7:0] mem_0_180_R0_data;
  wire  mem_0_180_R0_en;
  wire [6:0] mem_0_181_W0_addr;
  wire  mem_0_181_W0_clk;
  wire [7:0] mem_0_181_W0_data;
  wire  mem_0_181_W0_en;
  wire  mem_0_181_W0_mask;
  wire [6:0] mem_0_181_R0_addr;
  wire  mem_0_181_R0_clk;
  wire [7:0] mem_0_181_R0_data;
  wire  mem_0_181_R0_en;
  wire [6:0] mem_0_182_W0_addr;
  wire  mem_0_182_W0_clk;
  wire [7:0] mem_0_182_W0_data;
  wire  mem_0_182_W0_en;
  wire  mem_0_182_W0_mask;
  wire [6:0] mem_0_182_R0_addr;
  wire  mem_0_182_R0_clk;
  wire [7:0] mem_0_182_R0_data;
  wire  mem_0_182_R0_en;
  wire [6:0] mem_0_183_W0_addr;
  wire  mem_0_183_W0_clk;
  wire [7:0] mem_0_183_W0_data;
  wire  mem_0_183_W0_en;
  wire  mem_0_183_W0_mask;
  wire [6:0] mem_0_183_R0_addr;
  wire  mem_0_183_R0_clk;
  wire [7:0] mem_0_183_R0_data;
  wire  mem_0_183_R0_en;
  wire [6:0] mem_0_184_W0_addr;
  wire  mem_0_184_W0_clk;
  wire [7:0] mem_0_184_W0_data;
  wire  mem_0_184_W0_en;
  wire  mem_0_184_W0_mask;
  wire [6:0] mem_0_184_R0_addr;
  wire  mem_0_184_R0_clk;
  wire [7:0] mem_0_184_R0_data;
  wire  mem_0_184_R0_en;
  wire [6:0] mem_0_185_W0_addr;
  wire  mem_0_185_W0_clk;
  wire [7:0] mem_0_185_W0_data;
  wire  mem_0_185_W0_en;
  wire  mem_0_185_W0_mask;
  wire [6:0] mem_0_185_R0_addr;
  wire  mem_0_185_R0_clk;
  wire [7:0] mem_0_185_R0_data;
  wire  mem_0_185_R0_en;
  wire [6:0] mem_0_186_W0_addr;
  wire  mem_0_186_W0_clk;
  wire [7:0] mem_0_186_W0_data;
  wire  mem_0_186_W0_en;
  wire  mem_0_186_W0_mask;
  wire [6:0] mem_0_186_R0_addr;
  wire  mem_0_186_R0_clk;
  wire [7:0] mem_0_186_R0_data;
  wire  mem_0_186_R0_en;
  wire [6:0] mem_0_187_W0_addr;
  wire  mem_0_187_W0_clk;
  wire [7:0] mem_0_187_W0_data;
  wire  mem_0_187_W0_en;
  wire  mem_0_187_W0_mask;
  wire [6:0] mem_0_187_R0_addr;
  wire  mem_0_187_R0_clk;
  wire [7:0] mem_0_187_R0_data;
  wire  mem_0_187_R0_en;
  wire [6:0] mem_0_188_W0_addr;
  wire  mem_0_188_W0_clk;
  wire [7:0] mem_0_188_W0_data;
  wire  mem_0_188_W0_en;
  wire  mem_0_188_W0_mask;
  wire [6:0] mem_0_188_R0_addr;
  wire  mem_0_188_R0_clk;
  wire [7:0] mem_0_188_R0_data;
  wire  mem_0_188_R0_en;
  wire [6:0] mem_0_189_W0_addr;
  wire  mem_0_189_W0_clk;
  wire [7:0] mem_0_189_W0_data;
  wire  mem_0_189_W0_en;
  wire  mem_0_189_W0_mask;
  wire [6:0] mem_0_189_R0_addr;
  wire  mem_0_189_R0_clk;
  wire [7:0] mem_0_189_R0_data;
  wire  mem_0_189_R0_en;
  wire [6:0] mem_0_190_W0_addr;
  wire  mem_0_190_W0_clk;
  wire [7:0] mem_0_190_W0_data;
  wire  mem_0_190_W0_en;
  wire  mem_0_190_W0_mask;
  wire [6:0] mem_0_190_R0_addr;
  wire  mem_0_190_R0_clk;
  wire [7:0] mem_0_190_R0_data;
  wire  mem_0_190_R0_en;
  wire [6:0] mem_0_191_W0_addr;
  wire  mem_0_191_W0_clk;
  wire [7:0] mem_0_191_W0_data;
  wire  mem_0_191_W0_en;
  wire  mem_0_191_W0_mask;
  wire [6:0] mem_0_191_R0_addr;
  wire  mem_0_191_R0_clk;
  wire [7:0] mem_0_191_R0_data;
  wire  mem_0_191_R0_en;
  wire [6:0] mem_0_192_W0_addr;
  wire  mem_0_192_W0_clk;
  wire [7:0] mem_0_192_W0_data;
  wire  mem_0_192_W0_en;
  wire  mem_0_192_W0_mask;
  wire [6:0] mem_0_192_R0_addr;
  wire  mem_0_192_R0_clk;
  wire [7:0] mem_0_192_R0_data;
  wire  mem_0_192_R0_en;
  wire [6:0] mem_0_193_W0_addr;
  wire  mem_0_193_W0_clk;
  wire [7:0] mem_0_193_W0_data;
  wire  mem_0_193_W0_en;
  wire  mem_0_193_W0_mask;
  wire [6:0] mem_0_193_R0_addr;
  wire  mem_0_193_R0_clk;
  wire [7:0] mem_0_193_R0_data;
  wire  mem_0_193_R0_en;
  wire [6:0] mem_0_194_W0_addr;
  wire  mem_0_194_W0_clk;
  wire [7:0] mem_0_194_W0_data;
  wire  mem_0_194_W0_en;
  wire  mem_0_194_W0_mask;
  wire [6:0] mem_0_194_R0_addr;
  wire  mem_0_194_R0_clk;
  wire [7:0] mem_0_194_R0_data;
  wire  mem_0_194_R0_en;
  wire [6:0] mem_0_195_W0_addr;
  wire  mem_0_195_W0_clk;
  wire [7:0] mem_0_195_W0_data;
  wire  mem_0_195_W0_en;
  wire  mem_0_195_W0_mask;
  wire [6:0] mem_0_195_R0_addr;
  wire  mem_0_195_R0_clk;
  wire [7:0] mem_0_195_R0_data;
  wire  mem_0_195_R0_en;
  wire [6:0] mem_0_196_W0_addr;
  wire  mem_0_196_W0_clk;
  wire [7:0] mem_0_196_W0_data;
  wire  mem_0_196_W0_en;
  wire  mem_0_196_W0_mask;
  wire [6:0] mem_0_196_R0_addr;
  wire  mem_0_196_R0_clk;
  wire [7:0] mem_0_196_R0_data;
  wire  mem_0_196_R0_en;
  wire [6:0] mem_0_197_W0_addr;
  wire  mem_0_197_W0_clk;
  wire [7:0] mem_0_197_W0_data;
  wire  mem_0_197_W0_en;
  wire  mem_0_197_W0_mask;
  wire [6:0] mem_0_197_R0_addr;
  wire  mem_0_197_R0_clk;
  wire [7:0] mem_0_197_R0_data;
  wire  mem_0_197_R0_en;
  wire [6:0] mem_0_198_W0_addr;
  wire  mem_0_198_W0_clk;
  wire [7:0] mem_0_198_W0_data;
  wire  mem_0_198_W0_en;
  wire  mem_0_198_W0_mask;
  wire [6:0] mem_0_198_R0_addr;
  wire  mem_0_198_R0_clk;
  wire [7:0] mem_0_198_R0_data;
  wire  mem_0_198_R0_en;
  wire [6:0] mem_0_199_W0_addr;
  wire  mem_0_199_W0_clk;
  wire [7:0] mem_0_199_W0_data;
  wire  mem_0_199_W0_en;
  wire  mem_0_199_W0_mask;
  wire [6:0] mem_0_199_R0_addr;
  wire  mem_0_199_R0_clk;
  wire [7:0] mem_0_199_R0_data;
  wire  mem_0_199_R0_en;
  wire [6:0] mem_0_200_W0_addr;
  wire  mem_0_200_W0_clk;
  wire [7:0] mem_0_200_W0_data;
  wire  mem_0_200_W0_en;
  wire  mem_0_200_W0_mask;
  wire [6:0] mem_0_200_R0_addr;
  wire  mem_0_200_R0_clk;
  wire [7:0] mem_0_200_R0_data;
  wire  mem_0_200_R0_en;
  wire [6:0] mem_0_201_W0_addr;
  wire  mem_0_201_W0_clk;
  wire [7:0] mem_0_201_W0_data;
  wire  mem_0_201_W0_en;
  wire  mem_0_201_W0_mask;
  wire [6:0] mem_0_201_R0_addr;
  wire  mem_0_201_R0_clk;
  wire [7:0] mem_0_201_R0_data;
  wire  mem_0_201_R0_en;
  wire [6:0] mem_0_202_W0_addr;
  wire  mem_0_202_W0_clk;
  wire [7:0] mem_0_202_W0_data;
  wire  mem_0_202_W0_en;
  wire  mem_0_202_W0_mask;
  wire [6:0] mem_0_202_R0_addr;
  wire  mem_0_202_R0_clk;
  wire [7:0] mem_0_202_R0_data;
  wire  mem_0_202_R0_en;
  wire [6:0] mem_0_203_W0_addr;
  wire  mem_0_203_W0_clk;
  wire [7:0] mem_0_203_W0_data;
  wire  mem_0_203_W0_en;
  wire  mem_0_203_W0_mask;
  wire [6:0] mem_0_203_R0_addr;
  wire  mem_0_203_R0_clk;
  wire [7:0] mem_0_203_R0_data;
  wire  mem_0_203_R0_en;
  wire [6:0] mem_0_204_W0_addr;
  wire  mem_0_204_W0_clk;
  wire [7:0] mem_0_204_W0_data;
  wire  mem_0_204_W0_en;
  wire  mem_0_204_W0_mask;
  wire [6:0] mem_0_204_R0_addr;
  wire  mem_0_204_R0_clk;
  wire [7:0] mem_0_204_R0_data;
  wire  mem_0_204_R0_en;
  wire [6:0] mem_0_205_W0_addr;
  wire  mem_0_205_W0_clk;
  wire [7:0] mem_0_205_W0_data;
  wire  mem_0_205_W0_en;
  wire  mem_0_205_W0_mask;
  wire [6:0] mem_0_205_R0_addr;
  wire  mem_0_205_R0_clk;
  wire [7:0] mem_0_205_R0_data;
  wire  mem_0_205_R0_en;
  wire [6:0] mem_0_206_W0_addr;
  wire  mem_0_206_W0_clk;
  wire [7:0] mem_0_206_W0_data;
  wire  mem_0_206_W0_en;
  wire  mem_0_206_W0_mask;
  wire [6:0] mem_0_206_R0_addr;
  wire  mem_0_206_R0_clk;
  wire [7:0] mem_0_206_R0_data;
  wire  mem_0_206_R0_en;
  wire [6:0] mem_0_207_W0_addr;
  wire  mem_0_207_W0_clk;
  wire [7:0] mem_0_207_W0_data;
  wire  mem_0_207_W0_en;
  wire  mem_0_207_W0_mask;
  wire [6:0] mem_0_207_R0_addr;
  wire  mem_0_207_R0_clk;
  wire [7:0] mem_0_207_R0_data;
  wire  mem_0_207_R0_en;
  wire [6:0] mem_0_208_W0_addr;
  wire  mem_0_208_W0_clk;
  wire [7:0] mem_0_208_W0_data;
  wire  mem_0_208_W0_en;
  wire  mem_0_208_W0_mask;
  wire [6:0] mem_0_208_R0_addr;
  wire  mem_0_208_R0_clk;
  wire [7:0] mem_0_208_R0_data;
  wire  mem_0_208_R0_en;
  wire [6:0] mem_0_209_W0_addr;
  wire  mem_0_209_W0_clk;
  wire [7:0] mem_0_209_W0_data;
  wire  mem_0_209_W0_en;
  wire  mem_0_209_W0_mask;
  wire [6:0] mem_0_209_R0_addr;
  wire  mem_0_209_R0_clk;
  wire [7:0] mem_0_209_R0_data;
  wire  mem_0_209_R0_en;
  wire [6:0] mem_0_210_W0_addr;
  wire  mem_0_210_W0_clk;
  wire [7:0] mem_0_210_W0_data;
  wire  mem_0_210_W0_en;
  wire  mem_0_210_W0_mask;
  wire [6:0] mem_0_210_R0_addr;
  wire  mem_0_210_R0_clk;
  wire [7:0] mem_0_210_R0_data;
  wire  mem_0_210_R0_en;
  wire [6:0] mem_0_211_W0_addr;
  wire  mem_0_211_W0_clk;
  wire [7:0] mem_0_211_W0_data;
  wire  mem_0_211_W0_en;
  wire  mem_0_211_W0_mask;
  wire [6:0] mem_0_211_R0_addr;
  wire  mem_0_211_R0_clk;
  wire [7:0] mem_0_211_R0_data;
  wire  mem_0_211_R0_en;
  wire [6:0] mem_0_212_W0_addr;
  wire  mem_0_212_W0_clk;
  wire [7:0] mem_0_212_W0_data;
  wire  mem_0_212_W0_en;
  wire  mem_0_212_W0_mask;
  wire [6:0] mem_0_212_R0_addr;
  wire  mem_0_212_R0_clk;
  wire [7:0] mem_0_212_R0_data;
  wire  mem_0_212_R0_en;
  wire [6:0] mem_0_213_W0_addr;
  wire  mem_0_213_W0_clk;
  wire [7:0] mem_0_213_W0_data;
  wire  mem_0_213_W0_en;
  wire  mem_0_213_W0_mask;
  wire [6:0] mem_0_213_R0_addr;
  wire  mem_0_213_R0_clk;
  wire [7:0] mem_0_213_R0_data;
  wire  mem_0_213_R0_en;
  wire [6:0] mem_0_214_W0_addr;
  wire  mem_0_214_W0_clk;
  wire [7:0] mem_0_214_W0_data;
  wire  mem_0_214_W0_en;
  wire  mem_0_214_W0_mask;
  wire [6:0] mem_0_214_R0_addr;
  wire  mem_0_214_R0_clk;
  wire [7:0] mem_0_214_R0_data;
  wire  mem_0_214_R0_en;
  wire [6:0] mem_0_215_W0_addr;
  wire  mem_0_215_W0_clk;
  wire [7:0] mem_0_215_W0_data;
  wire  mem_0_215_W0_en;
  wire  mem_0_215_W0_mask;
  wire [6:0] mem_0_215_R0_addr;
  wire  mem_0_215_R0_clk;
  wire [7:0] mem_0_215_R0_data;
  wire  mem_0_215_R0_en;
  wire [6:0] mem_0_216_W0_addr;
  wire  mem_0_216_W0_clk;
  wire [7:0] mem_0_216_W0_data;
  wire  mem_0_216_W0_en;
  wire  mem_0_216_W0_mask;
  wire [6:0] mem_0_216_R0_addr;
  wire  mem_0_216_R0_clk;
  wire [7:0] mem_0_216_R0_data;
  wire  mem_0_216_R0_en;
  wire [6:0] mem_0_217_W0_addr;
  wire  mem_0_217_W0_clk;
  wire [7:0] mem_0_217_W0_data;
  wire  mem_0_217_W0_en;
  wire  mem_0_217_W0_mask;
  wire [6:0] mem_0_217_R0_addr;
  wire  mem_0_217_R0_clk;
  wire [7:0] mem_0_217_R0_data;
  wire  mem_0_217_R0_en;
  wire [6:0] mem_0_218_W0_addr;
  wire  mem_0_218_W0_clk;
  wire [7:0] mem_0_218_W0_data;
  wire  mem_0_218_W0_en;
  wire  mem_0_218_W0_mask;
  wire [6:0] mem_0_218_R0_addr;
  wire  mem_0_218_R0_clk;
  wire [7:0] mem_0_218_R0_data;
  wire  mem_0_218_R0_en;
  wire [6:0] mem_0_219_W0_addr;
  wire  mem_0_219_W0_clk;
  wire [7:0] mem_0_219_W0_data;
  wire  mem_0_219_W0_en;
  wire  mem_0_219_W0_mask;
  wire [6:0] mem_0_219_R0_addr;
  wire  mem_0_219_R0_clk;
  wire [7:0] mem_0_219_R0_data;
  wire  mem_0_219_R0_en;
  wire [6:0] mem_0_220_W0_addr;
  wire  mem_0_220_W0_clk;
  wire [7:0] mem_0_220_W0_data;
  wire  mem_0_220_W0_en;
  wire  mem_0_220_W0_mask;
  wire [6:0] mem_0_220_R0_addr;
  wire  mem_0_220_R0_clk;
  wire [7:0] mem_0_220_R0_data;
  wire  mem_0_220_R0_en;
  wire [6:0] mem_0_221_W0_addr;
  wire  mem_0_221_W0_clk;
  wire [7:0] mem_0_221_W0_data;
  wire  mem_0_221_W0_en;
  wire  mem_0_221_W0_mask;
  wire [6:0] mem_0_221_R0_addr;
  wire  mem_0_221_R0_clk;
  wire [7:0] mem_0_221_R0_data;
  wire  mem_0_221_R0_en;
  wire [6:0] mem_0_222_W0_addr;
  wire  mem_0_222_W0_clk;
  wire [7:0] mem_0_222_W0_data;
  wire  mem_0_222_W0_en;
  wire  mem_0_222_W0_mask;
  wire [6:0] mem_0_222_R0_addr;
  wire  mem_0_222_R0_clk;
  wire [7:0] mem_0_222_R0_data;
  wire  mem_0_222_R0_en;
  wire [6:0] mem_0_223_W0_addr;
  wire  mem_0_223_W0_clk;
  wire [7:0] mem_0_223_W0_data;
  wire  mem_0_223_W0_en;
  wire  mem_0_223_W0_mask;
  wire [6:0] mem_0_223_R0_addr;
  wire  mem_0_223_R0_clk;
  wire [7:0] mem_0_223_R0_data;
  wire  mem_0_223_R0_en;
  wire [6:0] mem_0_224_W0_addr;
  wire  mem_0_224_W0_clk;
  wire [7:0] mem_0_224_W0_data;
  wire  mem_0_224_W0_en;
  wire  mem_0_224_W0_mask;
  wire [6:0] mem_0_224_R0_addr;
  wire  mem_0_224_R0_clk;
  wire [7:0] mem_0_224_R0_data;
  wire  mem_0_224_R0_en;
  wire [6:0] mem_0_225_W0_addr;
  wire  mem_0_225_W0_clk;
  wire [7:0] mem_0_225_W0_data;
  wire  mem_0_225_W0_en;
  wire  mem_0_225_W0_mask;
  wire [6:0] mem_0_225_R0_addr;
  wire  mem_0_225_R0_clk;
  wire [7:0] mem_0_225_R0_data;
  wire  mem_0_225_R0_en;
  wire [6:0] mem_0_226_W0_addr;
  wire  mem_0_226_W0_clk;
  wire [7:0] mem_0_226_W0_data;
  wire  mem_0_226_W0_en;
  wire  mem_0_226_W0_mask;
  wire [6:0] mem_0_226_R0_addr;
  wire  mem_0_226_R0_clk;
  wire [7:0] mem_0_226_R0_data;
  wire  mem_0_226_R0_en;
  wire [6:0] mem_0_227_W0_addr;
  wire  mem_0_227_W0_clk;
  wire [7:0] mem_0_227_W0_data;
  wire  mem_0_227_W0_en;
  wire  mem_0_227_W0_mask;
  wire [6:0] mem_0_227_R0_addr;
  wire  mem_0_227_R0_clk;
  wire [7:0] mem_0_227_R0_data;
  wire  mem_0_227_R0_en;
  wire [6:0] mem_0_228_W0_addr;
  wire  mem_0_228_W0_clk;
  wire [7:0] mem_0_228_W0_data;
  wire  mem_0_228_W0_en;
  wire  mem_0_228_W0_mask;
  wire [6:0] mem_0_228_R0_addr;
  wire  mem_0_228_R0_clk;
  wire [7:0] mem_0_228_R0_data;
  wire  mem_0_228_R0_en;
  wire [6:0] mem_0_229_W0_addr;
  wire  mem_0_229_W0_clk;
  wire [7:0] mem_0_229_W0_data;
  wire  mem_0_229_W0_en;
  wire  mem_0_229_W0_mask;
  wire [6:0] mem_0_229_R0_addr;
  wire  mem_0_229_R0_clk;
  wire [7:0] mem_0_229_R0_data;
  wire  mem_0_229_R0_en;
  wire [6:0] mem_0_230_W0_addr;
  wire  mem_0_230_W0_clk;
  wire [7:0] mem_0_230_W0_data;
  wire  mem_0_230_W0_en;
  wire  mem_0_230_W0_mask;
  wire [6:0] mem_0_230_R0_addr;
  wire  mem_0_230_R0_clk;
  wire [7:0] mem_0_230_R0_data;
  wire  mem_0_230_R0_en;
  wire [6:0] mem_0_231_W0_addr;
  wire  mem_0_231_W0_clk;
  wire [7:0] mem_0_231_W0_data;
  wire  mem_0_231_W0_en;
  wire  mem_0_231_W0_mask;
  wire [6:0] mem_0_231_R0_addr;
  wire  mem_0_231_R0_clk;
  wire [7:0] mem_0_231_R0_data;
  wire  mem_0_231_R0_en;
  wire [6:0] mem_0_232_W0_addr;
  wire  mem_0_232_W0_clk;
  wire [7:0] mem_0_232_W0_data;
  wire  mem_0_232_W0_en;
  wire  mem_0_232_W0_mask;
  wire [6:0] mem_0_232_R0_addr;
  wire  mem_0_232_R0_clk;
  wire [7:0] mem_0_232_R0_data;
  wire  mem_0_232_R0_en;
  wire [6:0] mem_0_233_W0_addr;
  wire  mem_0_233_W0_clk;
  wire [7:0] mem_0_233_W0_data;
  wire  mem_0_233_W0_en;
  wire  mem_0_233_W0_mask;
  wire [6:0] mem_0_233_R0_addr;
  wire  mem_0_233_R0_clk;
  wire [7:0] mem_0_233_R0_data;
  wire  mem_0_233_R0_en;
  wire [6:0] mem_0_234_W0_addr;
  wire  mem_0_234_W0_clk;
  wire [7:0] mem_0_234_W0_data;
  wire  mem_0_234_W0_en;
  wire  mem_0_234_W0_mask;
  wire [6:0] mem_0_234_R0_addr;
  wire  mem_0_234_R0_clk;
  wire [7:0] mem_0_234_R0_data;
  wire  mem_0_234_R0_en;
  wire [6:0] mem_0_235_W0_addr;
  wire  mem_0_235_W0_clk;
  wire [7:0] mem_0_235_W0_data;
  wire  mem_0_235_W0_en;
  wire  mem_0_235_W0_mask;
  wire [6:0] mem_0_235_R0_addr;
  wire  mem_0_235_R0_clk;
  wire [7:0] mem_0_235_R0_data;
  wire  mem_0_235_R0_en;
  wire [6:0] mem_0_236_W0_addr;
  wire  mem_0_236_W0_clk;
  wire [7:0] mem_0_236_W0_data;
  wire  mem_0_236_W0_en;
  wire  mem_0_236_W0_mask;
  wire [6:0] mem_0_236_R0_addr;
  wire  mem_0_236_R0_clk;
  wire [7:0] mem_0_236_R0_data;
  wire  mem_0_236_R0_en;
  wire [6:0] mem_0_237_W0_addr;
  wire  mem_0_237_W0_clk;
  wire [7:0] mem_0_237_W0_data;
  wire  mem_0_237_W0_en;
  wire  mem_0_237_W0_mask;
  wire [6:0] mem_0_237_R0_addr;
  wire  mem_0_237_R0_clk;
  wire [7:0] mem_0_237_R0_data;
  wire  mem_0_237_R0_en;
  wire [6:0] mem_0_238_W0_addr;
  wire  mem_0_238_W0_clk;
  wire [7:0] mem_0_238_W0_data;
  wire  mem_0_238_W0_en;
  wire  mem_0_238_W0_mask;
  wire [6:0] mem_0_238_R0_addr;
  wire  mem_0_238_R0_clk;
  wire [7:0] mem_0_238_R0_data;
  wire  mem_0_238_R0_en;
  wire [6:0] mem_0_239_W0_addr;
  wire  mem_0_239_W0_clk;
  wire [7:0] mem_0_239_W0_data;
  wire  mem_0_239_W0_en;
  wire  mem_0_239_W0_mask;
  wire [6:0] mem_0_239_R0_addr;
  wire  mem_0_239_R0_clk;
  wire [7:0] mem_0_239_R0_data;
  wire  mem_0_239_R0_en;
  wire [6:0] mem_0_240_W0_addr;
  wire  mem_0_240_W0_clk;
  wire [7:0] mem_0_240_W0_data;
  wire  mem_0_240_W0_en;
  wire  mem_0_240_W0_mask;
  wire [6:0] mem_0_240_R0_addr;
  wire  mem_0_240_R0_clk;
  wire [7:0] mem_0_240_R0_data;
  wire  mem_0_240_R0_en;
  wire [6:0] mem_0_241_W0_addr;
  wire  mem_0_241_W0_clk;
  wire [7:0] mem_0_241_W0_data;
  wire  mem_0_241_W0_en;
  wire  mem_0_241_W0_mask;
  wire [6:0] mem_0_241_R0_addr;
  wire  mem_0_241_R0_clk;
  wire [7:0] mem_0_241_R0_data;
  wire  mem_0_241_R0_en;
  wire [6:0] mem_0_242_W0_addr;
  wire  mem_0_242_W0_clk;
  wire [7:0] mem_0_242_W0_data;
  wire  mem_0_242_W0_en;
  wire  mem_0_242_W0_mask;
  wire [6:0] mem_0_242_R0_addr;
  wire  mem_0_242_R0_clk;
  wire [7:0] mem_0_242_R0_data;
  wire  mem_0_242_R0_en;
  wire [6:0] mem_0_243_W0_addr;
  wire  mem_0_243_W0_clk;
  wire [7:0] mem_0_243_W0_data;
  wire  mem_0_243_W0_en;
  wire  mem_0_243_W0_mask;
  wire [6:0] mem_0_243_R0_addr;
  wire  mem_0_243_R0_clk;
  wire [7:0] mem_0_243_R0_data;
  wire  mem_0_243_R0_en;
  wire [6:0] mem_0_244_W0_addr;
  wire  mem_0_244_W0_clk;
  wire [7:0] mem_0_244_W0_data;
  wire  mem_0_244_W0_en;
  wire  mem_0_244_W0_mask;
  wire [6:0] mem_0_244_R0_addr;
  wire  mem_0_244_R0_clk;
  wire [7:0] mem_0_244_R0_data;
  wire  mem_0_244_R0_en;
  wire [6:0] mem_0_245_W0_addr;
  wire  mem_0_245_W0_clk;
  wire [7:0] mem_0_245_W0_data;
  wire  mem_0_245_W0_en;
  wire  mem_0_245_W0_mask;
  wire [6:0] mem_0_245_R0_addr;
  wire  mem_0_245_R0_clk;
  wire [7:0] mem_0_245_R0_data;
  wire  mem_0_245_R0_en;
  wire [6:0] mem_0_246_W0_addr;
  wire  mem_0_246_W0_clk;
  wire [7:0] mem_0_246_W0_data;
  wire  mem_0_246_W0_en;
  wire  mem_0_246_W0_mask;
  wire [6:0] mem_0_246_R0_addr;
  wire  mem_0_246_R0_clk;
  wire [7:0] mem_0_246_R0_data;
  wire  mem_0_246_R0_en;
  wire [6:0] mem_0_247_W0_addr;
  wire  mem_0_247_W0_clk;
  wire [7:0] mem_0_247_W0_data;
  wire  mem_0_247_W0_en;
  wire  mem_0_247_W0_mask;
  wire [6:0] mem_0_247_R0_addr;
  wire  mem_0_247_R0_clk;
  wire [7:0] mem_0_247_R0_data;
  wire  mem_0_247_R0_en;
  wire [6:0] mem_0_248_W0_addr;
  wire  mem_0_248_W0_clk;
  wire [7:0] mem_0_248_W0_data;
  wire  mem_0_248_W0_en;
  wire  mem_0_248_W0_mask;
  wire [6:0] mem_0_248_R0_addr;
  wire  mem_0_248_R0_clk;
  wire [7:0] mem_0_248_R0_data;
  wire  mem_0_248_R0_en;
  wire [6:0] mem_0_249_W0_addr;
  wire  mem_0_249_W0_clk;
  wire [7:0] mem_0_249_W0_data;
  wire  mem_0_249_W0_en;
  wire  mem_0_249_W0_mask;
  wire [6:0] mem_0_249_R0_addr;
  wire  mem_0_249_R0_clk;
  wire [7:0] mem_0_249_R0_data;
  wire  mem_0_249_R0_en;
  wire [6:0] mem_0_250_W0_addr;
  wire  mem_0_250_W0_clk;
  wire [7:0] mem_0_250_W0_data;
  wire  mem_0_250_W0_en;
  wire  mem_0_250_W0_mask;
  wire [6:0] mem_0_250_R0_addr;
  wire  mem_0_250_R0_clk;
  wire [7:0] mem_0_250_R0_data;
  wire  mem_0_250_R0_en;
  wire [6:0] mem_0_251_W0_addr;
  wire  mem_0_251_W0_clk;
  wire [7:0] mem_0_251_W0_data;
  wire  mem_0_251_W0_en;
  wire  mem_0_251_W0_mask;
  wire [6:0] mem_0_251_R0_addr;
  wire  mem_0_251_R0_clk;
  wire [7:0] mem_0_251_R0_data;
  wire  mem_0_251_R0_en;
  wire [6:0] mem_0_252_W0_addr;
  wire  mem_0_252_W0_clk;
  wire [7:0] mem_0_252_W0_data;
  wire  mem_0_252_W0_en;
  wire  mem_0_252_W0_mask;
  wire [6:0] mem_0_252_R0_addr;
  wire  mem_0_252_R0_clk;
  wire [7:0] mem_0_252_R0_data;
  wire  mem_0_252_R0_en;
  wire [6:0] mem_0_253_W0_addr;
  wire  mem_0_253_W0_clk;
  wire [7:0] mem_0_253_W0_data;
  wire  mem_0_253_W0_en;
  wire  mem_0_253_W0_mask;
  wire [6:0] mem_0_253_R0_addr;
  wire  mem_0_253_R0_clk;
  wire [7:0] mem_0_253_R0_data;
  wire  mem_0_253_R0_en;
  wire [6:0] mem_0_254_W0_addr;
  wire  mem_0_254_W0_clk;
  wire [7:0] mem_0_254_W0_data;
  wire  mem_0_254_W0_en;
  wire  mem_0_254_W0_mask;
  wire [6:0] mem_0_254_R0_addr;
  wire  mem_0_254_R0_clk;
  wire [7:0] mem_0_254_R0_data;
  wire  mem_0_254_R0_en;
  wire [6:0] mem_0_255_W0_addr;
  wire  mem_0_255_W0_clk;
  wire [7:0] mem_0_255_W0_data;
  wire  mem_0_255_W0_en;
  wire  mem_0_255_W0_mask;
  wire [6:0] mem_0_255_R0_addr;
  wire  mem_0_255_R0_clk;
  wire [7:0] mem_0_255_R0_data;
  wire  mem_0_255_R0_en;
  wire [7:0] R0_data_0_0 = mem_0_0_R0_data;
  wire [7:0] R0_data_0_1 = mem_0_1_R0_data;
  wire [7:0] R0_data_0_2 = mem_0_2_R0_data;
  wire [7:0] R0_data_0_3 = mem_0_3_R0_data;
  wire [7:0] R0_data_0_4 = mem_0_4_R0_data;
  wire [7:0] R0_data_0_5 = mem_0_5_R0_data;
  wire [7:0] R0_data_0_6 = mem_0_6_R0_data;
  wire [7:0] R0_data_0_7 = mem_0_7_R0_data;
  wire [7:0] R0_data_0_8 = mem_0_8_R0_data;
  wire [7:0] R0_data_0_9 = mem_0_9_R0_data;
  wire [7:0] R0_data_0_10 = mem_0_10_R0_data;
  wire [7:0] R0_data_0_11 = mem_0_11_R0_data;
  wire [7:0] R0_data_0_12 = mem_0_12_R0_data;
  wire [7:0] R0_data_0_13 = mem_0_13_R0_data;
  wire [7:0] R0_data_0_14 = mem_0_14_R0_data;
  wire [7:0] R0_data_0_15 = mem_0_15_R0_data;
  wire [7:0] R0_data_0_16 = mem_0_16_R0_data;
  wire [7:0] R0_data_0_17 = mem_0_17_R0_data;
  wire [7:0] R0_data_0_18 = mem_0_18_R0_data;
  wire [7:0] R0_data_0_19 = mem_0_19_R0_data;
  wire [7:0] R0_data_0_20 = mem_0_20_R0_data;
  wire [7:0] R0_data_0_21 = mem_0_21_R0_data;
  wire [7:0] R0_data_0_22 = mem_0_22_R0_data;
  wire [7:0] R0_data_0_23 = mem_0_23_R0_data;
  wire [7:0] R0_data_0_24 = mem_0_24_R0_data;
  wire [7:0] R0_data_0_25 = mem_0_25_R0_data;
  wire [7:0] R0_data_0_26 = mem_0_26_R0_data;
  wire [7:0] R0_data_0_27 = mem_0_27_R0_data;
  wire [7:0] R0_data_0_28 = mem_0_28_R0_data;
  wire [7:0] R0_data_0_29 = mem_0_29_R0_data;
  wire [7:0] R0_data_0_30 = mem_0_30_R0_data;
  wire [7:0] R0_data_0_31 = mem_0_31_R0_data;
  wire [7:0] R0_data_0_32 = mem_0_32_R0_data;
  wire [7:0] R0_data_0_33 = mem_0_33_R0_data;
  wire [7:0] R0_data_0_34 = mem_0_34_R0_data;
  wire [7:0] R0_data_0_35 = mem_0_35_R0_data;
  wire [7:0] R0_data_0_36 = mem_0_36_R0_data;
  wire [7:0] R0_data_0_37 = mem_0_37_R0_data;
  wire [7:0] R0_data_0_38 = mem_0_38_R0_data;
  wire [7:0] R0_data_0_39 = mem_0_39_R0_data;
  wire [7:0] R0_data_0_40 = mem_0_40_R0_data;
  wire [7:0] R0_data_0_41 = mem_0_41_R0_data;
  wire [7:0] R0_data_0_42 = mem_0_42_R0_data;
  wire [7:0] R0_data_0_43 = mem_0_43_R0_data;
  wire [7:0] R0_data_0_44 = mem_0_44_R0_data;
  wire [7:0] R0_data_0_45 = mem_0_45_R0_data;
  wire [7:0] R0_data_0_46 = mem_0_46_R0_data;
  wire [7:0] R0_data_0_47 = mem_0_47_R0_data;
  wire [7:0] R0_data_0_48 = mem_0_48_R0_data;
  wire [7:0] R0_data_0_49 = mem_0_49_R0_data;
  wire [7:0] R0_data_0_50 = mem_0_50_R0_data;
  wire [7:0] R0_data_0_51 = mem_0_51_R0_data;
  wire [7:0] R0_data_0_52 = mem_0_52_R0_data;
  wire [7:0] R0_data_0_53 = mem_0_53_R0_data;
  wire [7:0] R0_data_0_54 = mem_0_54_R0_data;
  wire [7:0] R0_data_0_55 = mem_0_55_R0_data;
  wire [7:0] R0_data_0_56 = mem_0_56_R0_data;
  wire [7:0] R0_data_0_57 = mem_0_57_R0_data;
  wire [7:0] R0_data_0_58 = mem_0_58_R0_data;
  wire [7:0] R0_data_0_59 = mem_0_59_R0_data;
  wire [7:0] R0_data_0_60 = mem_0_60_R0_data;
  wire [7:0] R0_data_0_61 = mem_0_61_R0_data;
  wire [7:0] R0_data_0_62 = mem_0_62_R0_data;
  wire [7:0] R0_data_0_63 = mem_0_63_R0_data;
  wire [7:0] R0_data_0_64 = mem_0_64_R0_data;
  wire [7:0] R0_data_0_65 = mem_0_65_R0_data;
  wire [7:0] R0_data_0_66 = mem_0_66_R0_data;
  wire [7:0] R0_data_0_67 = mem_0_67_R0_data;
  wire [7:0] R0_data_0_68 = mem_0_68_R0_data;
  wire [7:0] R0_data_0_69 = mem_0_69_R0_data;
  wire [7:0] R0_data_0_70 = mem_0_70_R0_data;
  wire [7:0] R0_data_0_71 = mem_0_71_R0_data;
  wire [7:0] R0_data_0_72 = mem_0_72_R0_data;
  wire [7:0] R0_data_0_73 = mem_0_73_R0_data;
  wire [7:0] R0_data_0_74 = mem_0_74_R0_data;
  wire [7:0] R0_data_0_75 = mem_0_75_R0_data;
  wire [7:0] R0_data_0_76 = mem_0_76_R0_data;
  wire [7:0] R0_data_0_77 = mem_0_77_R0_data;
  wire [7:0] R0_data_0_78 = mem_0_78_R0_data;
  wire [7:0] R0_data_0_79 = mem_0_79_R0_data;
  wire [7:0] R0_data_0_80 = mem_0_80_R0_data;
  wire [7:0] R0_data_0_81 = mem_0_81_R0_data;
  wire [7:0] R0_data_0_82 = mem_0_82_R0_data;
  wire [7:0] R0_data_0_83 = mem_0_83_R0_data;
  wire [7:0] R0_data_0_84 = mem_0_84_R0_data;
  wire [7:0] R0_data_0_85 = mem_0_85_R0_data;
  wire [7:0] R0_data_0_86 = mem_0_86_R0_data;
  wire [7:0] R0_data_0_87 = mem_0_87_R0_data;
  wire [7:0] R0_data_0_88 = mem_0_88_R0_data;
  wire [7:0] R0_data_0_89 = mem_0_89_R0_data;
  wire [7:0] R0_data_0_90 = mem_0_90_R0_data;
  wire [7:0] R0_data_0_91 = mem_0_91_R0_data;
  wire [7:0] R0_data_0_92 = mem_0_92_R0_data;
  wire [7:0] R0_data_0_93 = mem_0_93_R0_data;
  wire [7:0] R0_data_0_94 = mem_0_94_R0_data;
  wire [7:0] R0_data_0_95 = mem_0_95_R0_data;
  wire [7:0] R0_data_0_96 = mem_0_96_R0_data;
  wire [7:0] R0_data_0_97 = mem_0_97_R0_data;
  wire [7:0] R0_data_0_98 = mem_0_98_R0_data;
  wire [7:0] R0_data_0_99 = mem_0_99_R0_data;
  wire [7:0] R0_data_0_100 = mem_0_100_R0_data;
  wire [7:0] R0_data_0_101 = mem_0_101_R0_data;
  wire [7:0] R0_data_0_102 = mem_0_102_R0_data;
  wire [7:0] R0_data_0_103 = mem_0_103_R0_data;
  wire [7:0] R0_data_0_104 = mem_0_104_R0_data;
  wire [7:0] R0_data_0_105 = mem_0_105_R0_data;
  wire [7:0] R0_data_0_106 = mem_0_106_R0_data;
  wire [7:0] R0_data_0_107 = mem_0_107_R0_data;
  wire [7:0] R0_data_0_108 = mem_0_108_R0_data;
  wire [7:0] R0_data_0_109 = mem_0_109_R0_data;
  wire [7:0] R0_data_0_110 = mem_0_110_R0_data;
  wire [7:0] R0_data_0_111 = mem_0_111_R0_data;
  wire [7:0] R0_data_0_112 = mem_0_112_R0_data;
  wire [7:0] R0_data_0_113 = mem_0_113_R0_data;
  wire [7:0] R0_data_0_114 = mem_0_114_R0_data;
  wire [7:0] R0_data_0_115 = mem_0_115_R0_data;
  wire [7:0] R0_data_0_116 = mem_0_116_R0_data;
  wire [7:0] R0_data_0_117 = mem_0_117_R0_data;
  wire [7:0] R0_data_0_118 = mem_0_118_R0_data;
  wire [7:0] R0_data_0_119 = mem_0_119_R0_data;
  wire [7:0] R0_data_0_120 = mem_0_120_R0_data;
  wire [7:0] R0_data_0_121 = mem_0_121_R0_data;
  wire [7:0] R0_data_0_122 = mem_0_122_R0_data;
  wire [7:0] R0_data_0_123 = mem_0_123_R0_data;
  wire [7:0] R0_data_0_124 = mem_0_124_R0_data;
  wire [7:0] R0_data_0_125 = mem_0_125_R0_data;
  wire [7:0] R0_data_0_126 = mem_0_126_R0_data;
  wire [7:0] R0_data_0_127 = mem_0_127_R0_data;
  wire [7:0] R0_data_0_128 = mem_0_128_R0_data;
  wire [7:0] R0_data_0_129 = mem_0_129_R0_data;
  wire [7:0] R0_data_0_130 = mem_0_130_R0_data;
  wire [7:0] R0_data_0_131 = mem_0_131_R0_data;
  wire [7:0] R0_data_0_132 = mem_0_132_R0_data;
  wire [7:0] R0_data_0_133 = mem_0_133_R0_data;
  wire [7:0] R0_data_0_134 = mem_0_134_R0_data;
  wire [7:0] R0_data_0_135 = mem_0_135_R0_data;
  wire [7:0] R0_data_0_136 = mem_0_136_R0_data;
  wire [7:0] R0_data_0_137 = mem_0_137_R0_data;
  wire [7:0] R0_data_0_138 = mem_0_138_R0_data;
  wire [7:0] R0_data_0_139 = mem_0_139_R0_data;
  wire [7:0] R0_data_0_140 = mem_0_140_R0_data;
  wire [7:0] R0_data_0_141 = mem_0_141_R0_data;
  wire [7:0] R0_data_0_142 = mem_0_142_R0_data;
  wire [7:0] R0_data_0_143 = mem_0_143_R0_data;
  wire [7:0] R0_data_0_144 = mem_0_144_R0_data;
  wire [7:0] R0_data_0_145 = mem_0_145_R0_data;
  wire [7:0] R0_data_0_146 = mem_0_146_R0_data;
  wire [7:0] R0_data_0_147 = mem_0_147_R0_data;
  wire [7:0] R0_data_0_148 = mem_0_148_R0_data;
  wire [7:0] R0_data_0_149 = mem_0_149_R0_data;
  wire [7:0] R0_data_0_150 = mem_0_150_R0_data;
  wire [7:0] R0_data_0_151 = mem_0_151_R0_data;
  wire [7:0] R0_data_0_152 = mem_0_152_R0_data;
  wire [7:0] R0_data_0_153 = mem_0_153_R0_data;
  wire [7:0] R0_data_0_154 = mem_0_154_R0_data;
  wire [7:0] R0_data_0_155 = mem_0_155_R0_data;
  wire [7:0] R0_data_0_156 = mem_0_156_R0_data;
  wire [7:0] R0_data_0_157 = mem_0_157_R0_data;
  wire [7:0] R0_data_0_158 = mem_0_158_R0_data;
  wire [7:0] R0_data_0_159 = mem_0_159_R0_data;
  wire [7:0] R0_data_0_160 = mem_0_160_R0_data;
  wire [7:0] R0_data_0_161 = mem_0_161_R0_data;
  wire [7:0] R0_data_0_162 = mem_0_162_R0_data;
  wire [7:0] R0_data_0_163 = mem_0_163_R0_data;
  wire [7:0] R0_data_0_164 = mem_0_164_R0_data;
  wire [7:0] R0_data_0_165 = mem_0_165_R0_data;
  wire [7:0] R0_data_0_166 = mem_0_166_R0_data;
  wire [7:0] R0_data_0_167 = mem_0_167_R0_data;
  wire [7:0] R0_data_0_168 = mem_0_168_R0_data;
  wire [7:0] R0_data_0_169 = mem_0_169_R0_data;
  wire [7:0] R0_data_0_170 = mem_0_170_R0_data;
  wire [7:0] R0_data_0_171 = mem_0_171_R0_data;
  wire [7:0] R0_data_0_172 = mem_0_172_R0_data;
  wire [7:0] R0_data_0_173 = mem_0_173_R0_data;
  wire [7:0] R0_data_0_174 = mem_0_174_R0_data;
  wire [7:0] R0_data_0_175 = mem_0_175_R0_data;
  wire [7:0] R0_data_0_176 = mem_0_176_R0_data;
  wire [7:0] R0_data_0_177 = mem_0_177_R0_data;
  wire [7:0] R0_data_0_178 = mem_0_178_R0_data;
  wire [7:0] R0_data_0_179 = mem_0_179_R0_data;
  wire [7:0] R0_data_0_180 = mem_0_180_R0_data;
  wire [7:0] R0_data_0_181 = mem_0_181_R0_data;
  wire [7:0] R0_data_0_182 = mem_0_182_R0_data;
  wire [7:0] R0_data_0_183 = mem_0_183_R0_data;
  wire [7:0] R0_data_0_184 = mem_0_184_R0_data;
  wire [7:0] R0_data_0_185 = mem_0_185_R0_data;
  wire [7:0] R0_data_0_186 = mem_0_186_R0_data;
  wire [7:0] R0_data_0_187 = mem_0_187_R0_data;
  wire [7:0] R0_data_0_188 = mem_0_188_R0_data;
  wire [7:0] R0_data_0_189 = mem_0_189_R0_data;
  wire [7:0] R0_data_0_190 = mem_0_190_R0_data;
  wire [7:0] R0_data_0_191 = mem_0_191_R0_data;
  wire [7:0] R0_data_0_192 = mem_0_192_R0_data;
  wire [7:0] R0_data_0_193 = mem_0_193_R0_data;
  wire [7:0] R0_data_0_194 = mem_0_194_R0_data;
  wire [7:0] R0_data_0_195 = mem_0_195_R0_data;
  wire [7:0] R0_data_0_196 = mem_0_196_R0_data;
  wire [7:0] R0_data_0_197 = mem_0_197_R0_data;
  wire [7:0] R0_data_0_198 = mem_0_198_R0_data;
  wire [7:0] R0_data_0_199 = mem_0_199_R0_data;
  wire [7:0] R0_data_0_200 = mem_0_200_R0_data;
  wire [7:0] R0_data_0_201 = mem_0_201_R0_data;
  wire [7:0] R0_data_0_202 = mem_0_202_R0_data;
  wire [7:0] R0_data_0_203 = mem_0_203_R0_data;
  wire [7:0] R0_data_0_204 = mem_0_204_R0_data;
  wire [7:0] R0_data_0_205 = mem_0_205_R0_data;
  wire [7:0] R0_data_0_206 = mem_0_206_R0_data;
  wire [7:0] R0_data_0_207 = mem_0_207_R0_data;
  wire [7:0] R0_data_0_208 = mem_0_208_R0_data;
  wire [7:0] R0_data_0_209 = mem_0_209_R0_data;
  wire [7:0] R0_data_0_210 = mem_0_210_R0_data;
  wire [7:0] R0_data_0_211 = mem_0_211_R0_data;
  wire [7:0] R0_data_0_212 = mem_0_212_R0_data;
  wire [7:0] R0_data_0_213 = mem_0_213_R0_data;
  wire [7:0] R0_data_0_214 = mem_0_214_R0_data;
  wire [7:0] R0_data_0_215 = mem_0_215_R0_data;
  wire [7:0] R0_data_0_216 = mem_0_216_R0_data;
  wire [7:0] R0_data_0_217 = mem_0_217_R0_data;
  wire [7:0] R0_data_0_218 = mem_0_218_R0_data;
  wire [7:0] R0_data_0_219 = mem_0_219_R0_data;
  wire [7:0] R0_data_0_220 = mem_0_220_R0_data;
  wire [7:0] R0_data_0_221 = mem_0_221_R0_data;
  wire [7:0] R0_data_0_222 = mem_0_222_R0_data;
  wire [7:0] R0_data_0_223 = mem_0_223_R0_data;
  wire [7:0] R0_data_0_224 = mem_0_224_R0_data;
  wire [7:0] R0_data_0_225 = mem_0_225_R0_data;
  wire [7:0] R0_data_0_226 = mem_0_226_R0_data;
  wire [7:0] R0_data_0_227 = mem_0_227_R0_data;
  wire [7:0] R0_data_0_228 = mem_0_228_R0_data;
  wire [7:0] R0_data_0_229 = mem_0_229_R0_data;
  wire [7:0] R0_data_0_230 = mem_0_230_R0_data;
  wire [7:0] R0_data_0_231 = mem_0_231_R0_data;
  wire [7:0] R0_data_0_232 = mem_0_232_R0_data;
  wire [7:0] R0_data_0_233 = mem_0_233_R0_data;
  wire [7:0] R0_data_0_234 = mem_0_234_R0_data;
  wire [7:0] R0_data_0_235 = mem_0_235_R0_data;
  wire [7:0] R0_data_0_236 = mem_0_236_R0_data;
  wire [7:0] R0_data_0_237 = mem_0_237_R0_data;
  wire [7:0] R0_data_0_238 = mem_0_238_R0_data;
  wire [7:0] R0_data_0_239 = mem_0_239_R0_data;
  wire [7:0] R0_data_0_240 = mem_0_240_R0_data;
  wire [7:0] R0_data_0_241 = mem_0_241_R0_data;
  wire [7:0] R0_data_0_242 = mem_0_242_R0_data;
  wire [7:0] R0_data_0_243 = mem_0_243_R0_data;
  wire [7:0] R0_data_0_244 = mem_0_244_R0_data;
  wire [7:0] R0_data_0_245 = mem_0_245_R0_data;
  wire [7:0] R0_data_0_246 = mem_0_246_R0_data;
  wire [7:0] R0_data_0_247 = mem_0_247_R0_data;
  wire [7:0] R0_data_0_248 = mem_0_248_R0_data;
  wire [7:0] R0_data_0_249 = mem_0_249_R0_data;
  wire [7:0] R0_data_0_250 = mem_0_250_R0_data;
  wire [7:0] R0_data_0_251 = mem_0_251_R0_data;
  wire [7:0] R0_data_0_252 = mem_0_252_R0_data;
  wire [7:0] R0_data_0_253 = mem_0_253_R0_data;
  wire [7:0] R0_data_0_254 = mem_0_254_R0_data;
  wire [7:0] R0_data_0_255 = mem_0_255_R0_data;
  wire [15:0] _GEN_0 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_2 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_3 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_4 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_5 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_6 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}
    ;
  wire [71:0] _GEN_7 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,
    R0_data_0_0};
  wire [79:0] _GEN_8 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,
    R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_9 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_14 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_15 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_16 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_17 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_18 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_19 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_20 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_21 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_22 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_23 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_24 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_25 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_26 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_27 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_28 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_29 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_30 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_31 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_32 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_33 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_34 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_35 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_36 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_37 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_38 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_39 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_40 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_41 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_42 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_43 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_44 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_45 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_46 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_47 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_48 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_49 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_50 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_51 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_52 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_53 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_54 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_55 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_56 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_57 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_58 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_59 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_60 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_61 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  wire [511:0] _GEN_62 = {R0_data_0_63,R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,
    R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [519:0] _GEN_63 = {R0_data_0_64,_GEN_62};
  wire [527:0] _GEN_64 = {R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [535:0] _GEN_65 = {R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [543:0] _GEN_66 = {R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [551:0] _GEN_67 = {R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [559:0] _GEN_68 = {R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [567:0] _GEN_69 = {R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,
    _GEN_62};
  wire [575:0] _GEN_70 = {R0_data_0_71,R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,
    R0_data_0_64,_GEN_62};
  wire [583:0] _GEN_71 = {R0_data_0_72,R0_data_0_71,R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,
    R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [591:0] _GEN_72 = {R0_data_0_73,_GEN_71};
  wire [599:0] _GEN_73 = {R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [607:0] _GEN_74 = {R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [615:0] _GEN_75 = {R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [623:0] _GEN_76 = {R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [631:0] _GEN_77 = {R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [639:0] _GEN_78 = {R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,
    _GEN_71};
  wire [647:0] _GEN_79 = {R0_data_0_80,R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,
    R0_data_0_73,_GEN_71};
  wire [655:0] _GEN_80 = {R0_data_0_81,R0_data_0_80,R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,
    R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [663:0] _GEN_81 = {R0_data_0_82,_GEN_80};
  wire [671:0] _GEN_82 = {R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [679:0] _GEN_83 = {R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [687:0] _GEN_84 = {R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [695:0] _GEN_85 = {R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [703:0] _GEN_86 = {R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [711:0] _GEN_87 = {R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,
    _GEN_80};
  wire [719:0] _GEN_88 = {R0_data_0_89,R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,
    R0_data_0_82,_GEN_80};
  wire [727:0] _GEN_89 = {R0_data_0_90,R0_data_0_89,R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,
    R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [735:0] _GEN_90 = {R0_data_0_91,_GEN_89};
  wire [743:0] _GEN_91 = {R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [751:0] _GEN_92 = {R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [759:0] _GEN_93 = {R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [767:0] _GEN_94 = {R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [775:0] _GEN_95 = {R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [783:0] _GEN_96 = {R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,
    _GEN_89};
  wire [791:0] _GEN_97 = {R0_data_0_98,R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,
    R0_data_0_91,_GEN_89};
  wire [799:0] _GEN_98 = {R0_data_0_99,R0_data_0_98,R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,
    R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [807:0] _GEN_99 = {R0_data_0_100,_GEN_98};
  wire [815:0] _GEN_100 = {R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [823:0] _GEN_101 = {R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [831:0] _GEN_102 = {R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [839:0] _GEN_103 = {R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [847:0] _GEN_104 = {R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [855:0] _GEN_105 = {R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,
    R0_data_0_100,_GEN_98};
  wire [863:0] _GEN_106 = {R0_data_0_107,R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,
    R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [871:0] _GEN_107 = {R0_data_0_108,R0_data_0_107,R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,
    R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [879:0] _GEN_108 = {R0_data_0_109,_GEN_107};
  wire [887:0] _GEN_109 = {R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [895:0] _GEN_110 = {R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [903:0] _GEN_111 = {R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [911:0] _GEN_112 = {R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [919:0] _GEN_113 = {R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107}
    ;
  wire [927:0] _GEN_114 = {R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,
    R0_data_0_109,_GEN_107};
  wire [935:0] _GEN_115 = {R0_data_0_116,R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,
    R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [943:0] _GEN_116 = {R0_data_0_117,R0_data_0_116,R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,
    R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [951:0] _GEN_117 = {R0_data_0_118,_GEN_116};
  wire [959:0] _GEN_118 = {R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [967:0] _GEN_119 = {R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [975:0] _GEN_120 = {R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [983:0] _GEN_121 = {R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [991:0] _GEN_122 = {R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116}
    ;
  wire [999:0] _GEN_123 = {R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,
    R0_data_0_118,_GEN_116};
  wire [1007:0] _GEN_124 = {R0_data_0_125,R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,
    R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [1015:0] _GEN_125 = {R0_data_0_126,R0_data_0_125,R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,
    R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [1023:0] _GEN_126 = {R0_data_0_127,_GEN_125};
  wire [1031:0] _GEN_127 = {R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1039:0] _GEN_128 = {R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1047:0] _GEN_129 = {R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1055:0] _GEN_130 = {R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1063:0] _GEN_131 = {R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125
    };
  wire [1071:0] _GEN_132 = {R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,
    R0_data_0_127,_GEN_125};
  wire [1079:0] _GEN_133 = {R0_data_0_134,R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,
    R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1087:0] _GEN_134 = {R0_data_0_135,R0_data_0_134,R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,
    R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1095:0] _GEN_135 = {R0_data_0_136,_GEN_134};
  wire [1103:0] _GEN_136 = {R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1111:0] _GEN_137 = {R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1119:0] _GEN_138 = {R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1127:0] _GEN_139 = {R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1135:0] _GEN_140 = {R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134
    };
  wire [1143:0] _GEN_141 = {R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,
    R0_data_0_136,_GEN_134};
  wire [1151:0] _GEN_142 = {R0_data_0_143,R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,
    R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1159:0] _GEN_143 = {R0_data_0_144,R0_data_0_143,R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,
    R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1167:0] _GEN_144 = {R0_data_0_145,_GEN_143};
  wire [1175:0] _GEN_145 = {R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1183:0] _GEN_146 = {R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1191:0] _GEN_147 = {R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1199:0] _GEN_148 = {R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1207:0] _GEN_149 = {R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143
    };
  wire [1215:0] _GEN_150 = {R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,
    R0_data_0_145,_GEN_143};
  wire [1223:0] _GEN_151 = {R0_data_0_152,R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,
    R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1231:0] _GEN_152 = {R0_data_0_153,R0_data_0_152,R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,
    R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1239:0] _GEN_153 = {R0_data_0_154,_GEN_152};
  wire [1247:0] _GEN_154 = {R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1255:0] _GEN_155 = {R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1263:0] _GEN_156 = {R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1271:0] _GEN_157 = {R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1279:0] _GEN_158 = {R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152
    };
  wire [1287:0] _GEN_159 = {R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,
    R0_data_0_154,_GEN_152};
  wire [1295:0] _GEN_160 = {R0_data_0_161,R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,
    R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1303:0] _GEN_161 = {R0_data_0_162,R0_data_0_161,R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,
    R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1311:0] _GEN_162 = {R0_data_0_163,_GEN_161};
  wire [1319:0] _GEN_163 = {R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1327:0] _GEN_164 = {R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1335:0] _GEN_165 = {R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1343:0] _GEN_166 = {R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1351:0] _GEN_167 = {R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161
    };
  wire [1359:0] _GEN_168 = {R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,
    R0_data_0_163,_GEN_161};
  wire [1367:0] _GEN_169 = {R0_data_0_170,R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,
    R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1375:0] _GEN_170 = {R0_data_0_171,R0_data_0_170,R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,
    R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1383:0] _GEN_171 = {R0_data_0_172,_GEN_170};
  wire [1391:0] _GEN_172 = {R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1399:0] _GEN_173 = {R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1407:0] _GEN_174 = {R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1415:0] _GEN_175 = {R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1423:0] _GEN_176 = {R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170
    };
  wire [1431:0] _GEN_177 = {R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,
    R0_data_0_172,_GEN_170};
  wire [1439:0] _GEN_178 = {R0_data_0_179,R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,
    R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1447:0] _GEN_179 = {R0_data_0_180,R0_data_0_179,R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,
    R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1455:0] _GEN_180 = {R0_data_0_181,_GEN_179};
  wire [1463:0] _GEN_181 = {R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1471:0] _GEN_182 = {R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1479:0] _GEN_183 = {R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1487:0] _GEN_184 = {R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1495:0] _GEN_185 = {R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179
    };
  wire [1503:0] _GEN_186 = {R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,
    R0_data_0_181,_GEN_179};
  wire [1511:0] _GEN_187 = {R0_data_0_188,R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,
    R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1519:0] _GEN_188 = {R0_data_0_189,R0_data_0_188,R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,
    R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1527:0] _GEN_189 = {R0_data_0_190,_GEN_188};
  wire [1535:0] _GEN_190 = {R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1543:0] _GEN_191 = {R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1551:0] _GEN_192 = {R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1559:0] _GEN_193 = {R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1567:0] _GEN_194 = {R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188
    };
  wire [1575:0] _GEN_195 = {R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,
    R0_data_0_190,_GEN_188};
  wire [1583:0] _GEN_196 = {R0_data_0_197,R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,
    R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1591:0] _GEN_197 = {R0_data_0_198,R0_data_0_197,R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,
    R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1599:0] _GEN_198 = {R0_data_0_199,_GEN_197};
  wire [1607:0] _GEN_199 = {R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1615:0] _GEN_200 = {R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1623:0] _GEN_201 = {R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1631:0] _GEN_202 = {R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1639:0] _GEN_203 = {R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197
    };
  wire [1647:0] _GEN_204 = {R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,
    R0_data_0_199,_GEN_197};
  wire [1655:0] _GEN_205 = {R0_data_0_206,R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,
    R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1663:0] _GEN_206 = {R0_data_0_207,R0_data_0_206,R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,
    R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1671:0] _GEN_207 = {R0_data_0_208,_GEN_206};
  wire [1679:0] _GEN_208 = {R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1687:0] _GEN_209 = {R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1695:0] _GEN_210 = {R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1703:0] _GEN_211 = {R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1711:0] _GEN_212 = {R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206
    };
  wire [1719:0] _GEN_213 = {R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,
    R0_data_0_208,_GEN_206};
  wire [1727:0] _GEN_214 = {R0_data_0_215,R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,
    R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1735:0] _GEN_215 = {R0_data_0_216,R0_data_0_215,R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,
    R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1743:0] _GEN_216 = {R0_data_0_217,_GEN_215};
  wire [1751:0] _GEN_217 = {R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1759:0] _GEN_218 = {R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1767:0] _GEN_219 = {R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1775:0] _GEN_220 = {R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1783:0] _GEN_221 = {R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215
    };
  wire [1791:0] _GEN_222 = {R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,
    R0_data_0_217,_GEN_215};
  wire [1799:0] _GEN_223 = {R0_data_0_224,R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,
    R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1807:0] _GEN_224 = {R0_data_0_225,R0_data_0_224,R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,
    R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1815:0] _GEN_225 = {R0_data_0_226,_GEN_224};
  wire [1823:0] _GEN_226 = {R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1831:0] _GEN_227 = {R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1839:0] _GEN_228 = {R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1847:0] _GEN_229 = {R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1855:0] _GEN_230 = {R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224
    };
  wire [1863:0] _GEN_231 = {R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,
    R0_data_0_226,_GEN_224};
  wire [1871:0] _GEN_232 = {R0_data_0_233,R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,
    R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1879:0] _GEN_233 = {R0_data_0_234,R0_data_0_233,R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,
    R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1887:0] _GEN_234 = {R0_data_0_235,_GEN_233};
  wire [1895:0] _GEN_235 = {R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1903:0] _GEN_236 = {R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1911:0] _GEN_237 = {R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1919:0] _GEN_238 = {R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1927:0] _GEN_239 = {R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233
    };
  wire [1935:0] _GEN_240 = {R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,
    R0_data_0_235,_GEN_233};
  wire [1943:0] _GEN_241 = {R0_data_0_242,R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,
    R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1951:0] _GEN_242 = {R0_data_0_243,R0_data_0_242,R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,
    R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1959:0] _GEN_243 = {R0_data_0_244,_GEN_242};
  wire [1967:0] _GEN_244 = {R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1975:0] _GEN_245 = {R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1983:0] _GEN_246 = {R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1991:0] _GEN_247 = {R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1999:0] _GEN_248 = {R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242
    };
  wire [2007:0] _GEN_249 = {R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,
    R0_data_0_244,_GEN_242};
  wire [2015:0] _GEN_250 = {R0_data_0_251,R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,
    R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [2023:0] _GEN_251 = {R0_data_0_252,R0_data_0_251,R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,
    R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [2031:0] _GEN_252 = {R0_data_0_253,_GEN_251};
  wire [2039:0] _GEN_253 = {R0_data_0_254,R0_data_0_253,_GEN_251};
  wire [2047:0] R0_data_0 = {R0_data_0_255,R0_data_0_254,R0_data_0_253,_GEN_251};
  wire [15:0] _GEN_254 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_255 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_256 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_257 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_258 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_259 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_260 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,
    R0_data_0_0};
  wire [71:0] _GEN_261 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,
    R0_data_0_1,R0_data_0_0};
  wire [79:0] _GEN_262 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,
    R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_263 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_264 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_265 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_266 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_267 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_268 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_269 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_270 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_271 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_272 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_273 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_274 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_275 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_276 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_277 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_278 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_279 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_280 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_281 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_282 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_283 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_284 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_285 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_286 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_287 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_288 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_289 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_290 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_291 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_292 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_293 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_294 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_295 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_296 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_297 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_298 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_299 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_300 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_301 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_302 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_303 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_304 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_305 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_306 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_307 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_308 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_309 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_310 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_311 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_312 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_313 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_314 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_315 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  wire [511:0] _GEN_316 = {R0_data_0_63,R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,
    R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [519:0] _GEN_317 = {R0_data_0_64,_GEN_62};
  wire [527:0] _GEN_318 = {R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [535:0] _GEN_319 = {R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [543:0] _GEN_320 = {R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [551:0] _GEN_321 = {R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [559:0] _GEN_322 = {R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [567:0] _GEN_323 = {R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,R0_data_0_64,
    _GEN_62};
  wire [575:0] _GEN_324 = {R0_data_0_71,R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,R0_data_0_65,
    R0_data_0_64,_GEN_62};
  wire [583:0] _GEN_325 = {R0_data_0_72,R0_data_0_71,R0_data_0_70,R0_data_0_69,R0_data_0_68,R0_data_0_67,R0_data_0_66,
    R0_data_0_65,R0_data_0_64,_GEN_62};
  wire [591:0] _GEN_326 = {R0_data_0_73,_GEN_71};
  wire [599:0] _GEN_327 = {R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [607:0] _GEN_328 = {R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [615:0] _GEN_329 = {R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [623:0] _GEN_330 = {R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [631:0] _GEN_331 = {R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [639:0] _GEN_332 = {R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,R0_data_0_73,
    _GEN_71};
  wire [647:0] _GEN_333 = {R0_data_0_80,R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,R0_data_0_74,
    R0_data_0_73,_GEN_71};
  wire [655:0] _GEN_334 = {R0_data_0_81,R0_data_0_80,R0_data_0_79,R0_data_0_78,R0_data_0_77,R0_data_0_76,R0_data_0_75,
    R0_data_0_74,R0_data_0_73,_GEN_71};
  wire [663:0] _GEN_335 = {R0_data_0_82,_GEN_80};
  wire [671:0] _GEN_336 = {R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [679:0] _GEN_337 = {R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [687:0] _GEN_338 = {R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [695:0] _GEN_339 = {R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [703:0] _GEN_340 = {R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [711:0] _GEN_341 = {R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,R0_data_0_82,
    _GEN_80};
  wire [719:0] _GEN_342 = {R0_data_0_89,R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,R0_data_0_83,
    R0_data_0_82,_GEN_80};
  wire [727:0] _GEN_343 = {R0_data_0_90,R0_data_0_89,R0_data_0_88,R0_data_0_87,R0_data_0_86,R0_data_0_85,R0_data_0_84,
    R0_data_0_83,R0_data_0_82,_GEN_80};
  wire [735:0] _GEN_344 = {R0_data_0_91,_GEN_89};
  wire [743:0] _GEN_345 = {R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [751:0] _GEN_346 = {R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [759:0] _GEN_347 = {R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [767:0] _GEN_348 = {R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [775:0] _GEN_349 = {R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [783:0] _GEN_350 = {R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,R0_data_0_91,
    _GEN_89};
  wire [791:0] _GEN_351 = {R0_data_0_98,R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,R0_data_0_92,
    R0_data_0_91,_GEN_89};
  wire [799:0] _GEN_352 = {R0_data_0_99,R0_data_0_98,R0_data_0_97,R0_data_0_96,R0_data_0_95,R0_data_0_94,R0_data_0_93,
    R0_data_0_92,R0_data_0_91,_GEN_89};
  wire [807:0] _GEN_353 = {R0_data_0_100,_GEN_98};
  wire [815:0] _GEN_354 = {R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [823:0] _GEN_355 = {R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [831:0] _GEN_356 = {R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [839:0] _GEN_357 = {R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [847:0] _GEN_358 = {R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [855:0] _GEN_359 = {R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,R0_data_0_101,
    R0_data_0_100,_GEN_98};
  wire [863:0] _GEN_360 = {R0_data_0_107,R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,R0_data_0_102,
    R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [871:0] _GEN_361 = {R0_data_0_108,R0_data_0_107,R0_data_0_106,R0_data_0_105,R0_data_0_104,R0_data_0_103,
    R0_data_0_102,R0_data_0_101,R0_data_0_100,_GEN_98};
  wire [879:0] _GEN_362 = {R0_data_0_109,_GEN_107};
  wire [887:0] _GEN_363 = {R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [895:0] _GEN_364 = {R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [903:0] _GEN_365 = {R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [911:0] _GEN_366 = {R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [919:0] _GEN_367 = {R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107}
    ;
  wire [927:0] _GEN_368 = {R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,R0_data_0_110,
    R0_data_0_109,_GEN_107};
  wire [935:0] _GEN_369 = {R0_data_0_116,R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,R0_data_0_111,
    R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [943:0] _GEN_370 = {R0_data_0_117,R0_data_0_116,R0_data_0_115,R0_data_0_114,R0_data_0_113,R0_data_0_112,
    R0_data_0_111,R0_data_0_110,R0_data_0_109,_GEN_107};
  wire [951:0] _GEN_371 = {R0_data_0_118,_GEN_116};
  wire [959:0] _GEN_372 = {R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [967:0] _GEN_373 = {R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [975:0] _GEN_374 = {R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [983:0] _GEN_375 = {R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [991:0] _GEN_376 = {R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116}
    ;
  wire [999:0] _GEN_377 = {R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,R0_data_0_119,
    R0_data_0_118,_GEN_116};
  wire [1007:0] _GEN_378 = {R0_data_0_125,R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,R0_data_0_120,
    R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [1015:0] _GEN_379 = {R0_data_0_126,R0_data_0_125,R0_data_0_124,R0_data_0_123,R0_data_0_122,R0_data_0_121,
    R0_data_0_120,R0_data_0_119,R0_data_0_118,_GEN_116};
  wire [1023:0] _GEN_380 = {R0_data_0_127,_GEN_125};
  wire [1031:0] _GEN_381 = {R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1039:0] _GEN_382 = {R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1047:0] _GEN_383 = {R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1055:0] _GEN_384 = {R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1063:0] _GEN_385 = {R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125
    };
  wire [1071:0] _GEN_386 = {R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,R0_data_0_128,
    R0_data_0_127,_GEN_125};
  wire [1079:0] _GEN_387 = {R0_data_0_134,R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,R0_data_0_129,
    R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1087:0] _GEN_388 = {R0_data_0_135,R0_data_0_134,R0_data_0_133,R0_data_0_132,R0_data_0_131,R0_data_0_130,
    R0_data_0_129,R0_data_0_128,R0_data_0_127,_GEN_125};
  wire [1095:0] _GEN_389 = {R0_data_0_136,_GEN_134};
  wire [1103:0] _GEN_390 = {R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1111:0] _GEN_391 = {R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1119:0] _GEN_392 = {R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1127:0] _GEN_393 = {R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1135:0] _GEN_394 = {R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134
    };
  wire [1143:0] _GEN_395 = {R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,R0_data_0_137,
    R0_data_0_136,_GEN_134};
  wire [1151:0] _GEN_396 = {R0_data_0_143,R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,R0_data_0_138,
    R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1159:0] _GEN_397 = {R0_data_0_144,R0_data_0_143,R0_data_0_142,R0_data_0_141,R0_data_0_140,R0_data_0_139,
    R0_data_0_138,R0_data_0_137,R0_data_0_136,_GEN_134};
  wire [1167:0] _GEN_398 = {R0_data_0_145,_GEN_143};
  wire [1175:0] _GEN_399 = {R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1183:0] _GEN_400 = {R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1191:0] _GEN_401 = {R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1199:0] _GEN_402 = {R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1207:0] _GEN_403 = {R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143
    };
  wire [1215:0] _GEN_404 = {R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,R0_data_0_146,
    R0_data_0_145,_GEN_143};
  wire [1223:0] _GEN_405 = {R0_data_0_152,R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,R0_data_0_147,
    R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1231:0] _GEN_406 = {R0_data_0_153,R0_data_0_152,R0_data_0_151,R0_data_0_150,R0_data_0_149,R0_data_0_148,
    R0_data_0_147,R0_data_0_146,R0_data_0_145,_GEN_143};
  wire [1239:0] _GEN_407 = {R0_data_0_154,_GEN_152};
  wire [1247:0] _GEN_408 = {R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1255:0] _GEN_409 = {R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1263:0] _GEN_410 = {R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1271:0] _GEN_411 = {R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1279:0] _GEN_412 = {R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152
    };
  wire [1287:0] _GEN_413 = {R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,R0_data_0_155,
    R0_data_0_154,_GEN_152};
  wire [1295:0] _GEN_414 = {R0_data_0_161,R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,R0_data_0_156,
    R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1303:0] _GEN_415 = {R0_data_0_162,R0_data_0_161,R0_data_0_160,R0_data_0_159,R0_data_0_158,R0_data_0_157,
    R0_data_0_156,R0_data_0_155,R0_data_0_154,_GEN_152};
  wire [1311:0] _GEN_416 = {R0_data_0_163,_GEN_161};
  wire [1319:0] _GEN_417 = {R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1327:0] _GEN_418 = {R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1335:0] _GEN_419 = {R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1343:0] _GEN_420 = {R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1351:0] _GEN_421 = {R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161
    };
  wire [1359:0] _GEN_422 = {R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,R0_data_0_164,
    R0_data_0_163,_GEN_161};
  wire [1367:0] _GEN_423 = {R0_data_0_170,R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,R0_data_0_165,
    R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1375:0] _GEN_424 = {R0_data_0_171,R0_data_0_170,R0_data_0_169,R0_data_0_168,R0_data_0_167,R0_data_0_166,
    R0_data_0_165,R0_data_0_164,R0_data_0_163,_GEN_161};
  wire [1383:0] _GEN_425 = {R0_data_0_172,_GEN_170};
  wire [1391:0] _GEN_426 = {R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1399:0] _GEN_427 = {R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1407:0] _GEN_428 = {R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1415:0] _GEN_429 = {R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1423:0] _GEN_430 = {R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170
    };
  wire [1431:0] _GEN_431 = {R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,R0_data_0_173,
    R0_data_0_172,_GEN_170};
  wire [1439:0] _GEN_432 = {R0_data_0_179,R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,R0_data_0_174,
    R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1447:0] _GEN_433 = {R0_data_0_180,R0_data_0_179,R0_data_0_178,R0_data_0_177,R0_data_0_176,R0_data_0_175,
    R0_data_0_174,R0_data_0_173,R0_data_0_172,_GEN_170};
  wire [1455:0] _GEN_434 = {R0_data_0_181,_GEN_179};
  wire [1463:0] _GEN_435 = {R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1471:0] _GEN_436 = {R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1479:0] _GEN_437 = {R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1487:0] _GEN_438 = {R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1495:0] _GEN_439 = {R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179
    };
  wire [1503:0] _GEN_440 = {R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,R0_data_0_182,
    R0_data_0_181,_GEN_179};
  wire [1511:0] _GEN_441 = {R0_data_0_188,R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,R0_data_0_183,
    R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1519:0] _GEN_442 = {R0_data_0_189,R0_data_0_188,R0_data_0_187,R0_data_0_186,R0_data_0_185,R0_data_0_184,
    R0_data_0_183,R0_data_0_182,R0_data_0_181,_GEN_179};
  wire [1527:0] _GEN_443 = {R0_data_0_190,_GEN_188};
  wire [1535:0] _GEN_444 = {R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1543:0] _GEN_445 = {R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1551:0] _GEN_446 = {R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1559:0] _GEN_447 = {R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1567:0] _GEN_448 = {R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188
    };
  wire [1575:0] _GEN_449 = {R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,R0_data_0_191,
    R0_data_0_190,_GEN_188};
  wire [1583:0] _GEN_450 = {R0_data_0_197,R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,R0_data_0_192,
    R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1591:0] _GEN_451 = {R0_data_0_198,R0_data_0_197,R0_data_0_196,R0_data_0_195,R0_data_0_194,R0_data_0_193,
    R0_data_0_192,R0_data_0_191,R0_data_0_190,_GEN_188};
  wire [1599:0] _GEN_452 = {R0_data_0_199,_GEN_197};
  wire [1607:0] _GEN_453 = {R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1615:0] _GEN_454 = {R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1623:0] _GEN_455 = {R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1631:0] _GEN_456 = {R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1639:0] _GEN_457 = {R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197
    };
  wire [1647:0] _GEN_458 = {R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,R0_data_0_200,
    R0_data_0_199,_GEN_197};
  wire [1655:0] _GEN_459 = {R0_data_0_206,R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,R0_data_0_201,
    R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1663:0] _GEN_460 = {R0_data_0_207,R0_data_0_206,R0_data_0_205,R0_data_0_204,R0_data_0_203,R0_data_0_202,
    R0_data_0_201,R0_data_0_200,R0_data_0_199,_GEN_197};
  wire [1671:0] _GEN_461 = {R0_data_0_208,_GEN_206};
  wire [1679:0] _GEN_462 = {R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1687:0] _GEN_463 = {R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1695:0] _GEN_464 = {R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1703:0] _GEN_465 = {R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1711:0] _GEN_466 = {R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206
    };
  wire [1719:0] _GEN_467 = {R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,R0_data_0_209,
    R0_data_0_208,_GEN_206};
  wire [1727:0] _GEN_468 = {R0_data_0_215,R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,R0_data_0_210,
    R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1735:0] _GEN_469 = {R0_data_0_216,R0_data_0_215,R0_data_0_214,R0_data_0_213,R0_data_0_212,R0_data_0_211,
    R0_data_0_210,R0_data_0_209,R0_data_0_208,_GEN_206};
  wire [1743:0] _GEN_470 = {R0_data_0_217,_GEN_215};
  wire [1751:0] _GEN_471 = {R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1759:0] _GEN_472 = {R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1767:0] _GEN_473 = {R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1775:0] _GEN_474 = {R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1783:0] _GEN_475 = {R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215
    };
  wire [1791:0] _GEN_476 = {R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,R0_data_0_218,
    R0_data_0_217,_GEN_215};
  wire [1799:0] _GEN_477 = {R0_data_0_224,R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,R0_data_0_219,
    R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1807:0] _GEN_478 = {R0_data_0_225,R0_data_0_224,R0_data_0_223,R0_data_0_222,R0_data_0_221,R0_data_0_220,
    R0_data_0_219,R0_data_0_218,R0_data_0_217,_GEN_215};
  wire [1815:0] _GEN_479 = {R0_data_0_226,_GEN_224};
  wire [1823:0] _GEN_480 = {R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1831:0] _GEN_481 = {R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1839:0] _GEN_482 = {R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1847:0] _GEN_483 = {R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1855:0] _GEN_484 = {R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224
    };
  wire [1863:0] _GEN_485 = {R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,R0_data_0_227,
    R0_data_0_226,_GEN_224};
  wire [1871:0] _GEN_486 = {R0_data_0_233,R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,R0_data_0_228,
    R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1879:0] _GEN_487 = {R0_data_0_234,R0_data_0_233,R0_data_0_232,R0_data_0_231,R0_data_0_230,R0_data_0_229,
    R0_data_0_228,R0_data_0_227,R0_data_0_226,_GEN_224};
  wire [1887:0] _GEN_488 = {R0_data_0_235,_GEN_233};
  wire [1895:0] _GEN_489 = {R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1903:0] _GEN_490 = {R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1911:0] _GEN_491 = {R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1919:0] _GEN_492 = {R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1927:0] _GEN_493 = {R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233
    };
  wire [1935:0] _GEN_494 = {R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,R0_data_0_236,
    R0_data_0_235,_GEN_233};
  wire [1943:0] _GEN_495 = {R0_data_0_242,R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,R0_data_0_237,
    R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1951:0] _GEN_496 = {R0_data_0_243,R0_data_0_242,R0_data_0_241,R0_data_0_240,R0_data_0_239,R0_data_0_238,
    R0_data_0_237,R0_data_0_236,R0_data_0_235,_GEN_233};
  wire [1959:0] _GEN_497 = {R0_data_0_244,_GEN_242};
  wire [1967:0] _GEN_498 = {R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1975:0] _GEN_499 = {R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1983:0] _GEN_500 = {R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1991:0] _GEN_501 = {R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [1999:0] _GEN_502 = {R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242
    };
  wire [2007:0] _GEN_503 = {R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,R0_data_0_245,
    R0_data_0_244,_GEN_242};
  wire [2015:0] _GEN_504 = {R0_data_0_251,R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,R0_data_0_246,
    R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [2023:0] _GEN_505 = {R0_data_0_252,R0_data_0_251,R0_data_0_250,R0_data_0_249,R0_data_0_248,R0_data_0_247,
    R0_data_0_246,R0_data_0_245,R0_data_0_244,_GEN_242};
  wire [2031:0] _GEN_506 = {R0_data_0_253,_GEN_251};
  wire [2039:0] _GEN_507 = {R0_data_0_254,R0_data_0_253,_GEN_251};
  split_mem_0_ext mem_0_0 (
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_mem_0_ext mem_0_1 (
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_mem_0_ext mem_0_2 (
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_mem_0_ext mem_0_3 (
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  split_mem_0_ext mem_0_4 (
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask),
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en)
  );
  split_mem_0_ext mem_0_5 (
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask),
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en)
  );
  split_mem_0_ext mem_0_6 (
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask),
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en)
  );
  split_mem_0_ext mem_0_7 (
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask),
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en)
  );
  split_mem_0_ext mem_0_8 (
    .W0_addr(mem_0_8_W0_addr),
    .W0_clk(mem_0_8_W0_clk),
    .W0_data(mem_0_8_W0_data),
    .W0_en(mem_0_8_W0_en),
    .W0_mask(mem_0_8_W0_mask),
    .R0_addr(mem_0_8_R0_addr),
    .R0_clk(mem_0_8_R0_clk),
    .R0_data(mem_0_8_R0_data),
    .R0_en(mem_0_8_R0_en)
  );
  split_mem_0_ext mem_0_9 (
    .W0_addr(mem_0_9_W0_addr),
    .W0_clk(mem_0_9_W0_clk),
    .W0_data(mem_0_9_W0_data),
    .W0_en(mem_0_9_W0_en),
    .W0_mask(mem_0_9_W0_mask),
    .R0_addr(mem_0_9_R0_addr),
    .R0_clk(mem_0_9_R0_clk),
    .R0_data(mem_0_9_R0_data),
    .R0_en(mem_0_9_R0_en)
  );
  split_mem_0_ext mem_0_10 (
    .W0_addr(mem_0_10_W0_addr),
    .W0_clk(mem_0_10_W0_clk),
    .W0_data(mem_0_10_W0_data),
    .W0_en(mem_0_10_W0_en),
    .W0_mask(mem_0_10_W0_mask),
    .R0_addr(mem_0_10_R0_addr),
    .R0_clk(mem_0_10_R0_clk),
    .R0_data(mem_0_10_R0_data),
    .R0_en(mem_0_10_R0_en)
  );
  split_mem_0_ext mem_0_11 (
    .W0_addr(mem_0_11_W0_addr),
    .W0_clk(mem_0_11_W0_clk),
    .W0_data(mem_0_11_W0_data),
    .W0_en(mem_0_11_W0_en),
    .W0_mask(mem_0_11_W0_mask),
    .R0_addr(mem_0_11_R0_addr),
    .R0_clk(mem_0_11_R0_clk),
    .R0_data(mem_0_11_R0_data),
    .R0_en(mem_0_11_R0_en)
  );
  split_mem_0_ext mem_0_12 (
    .W0_addr(mem_0_12_W0_addr),
    .W0_clk(mem_0_12_W0_clk),
    .W0_data(mem_0_12_W0_data),
    .W0_en(mem_0_12_W0_en),
    .W0_mask(mem_0_12_W0_mask),
    .R0_addr(mem_0_12_R0_addr),
    .R0_clk(mem_0_12_R0_clk),
    .R0_data(mem_0_12_R0_data),
    .R0_en(mem_0_12_R0_en)
  );
  split_mem_0_ext mem_0_13 (
    .W0_addr(mem_0_13_W0_addr),
    .W0_clk(mem_0_13_W0_clk),
    .W0_data(mem_0_13_W0_data),
    .W0_en(mem_0_13_W0_en),
    .W0_mask(mem_0_13_W0_mask),
    .R0_addr(mem_0_13_R0_addr),
    .R0_clk(mem_0_13_R0_clk),
    .R0_data(mem_0_13_R0_data),
    .R0_en(mem_0_13_R0_en)
  );
  split_mem_0_ext mem_0_14 (
    .W0_addr(mem_0_14_W0_addr),
    .W0_clk(mem_0_14_W0_clk),
    .W0_data(mem_0_14_W0_data),
    .W0_en(mem_0_14_W0_en),
    .W0_mask(mem_0_14_W0_mask),
    .R0_addr(mem_0_14_R0_addr),
    .R0_clk(mem_0_14_R0_clk),
    .R0_data(mem_0_14_R0_data),
    .R0_en(mem_0_14_R0_en)
  );
  split_mem_0_ext mem_0_15 (
    .W0_addr(mem_0_15_W0_addr),
    .W0_clk(mem_0_15_W0_clk),
    .W0_data(mem_0_15_W0_data),
    .W0_en(mem_0_15_W0_en),
    .W0_mask(mem_0_15_W0_mask),
    .R0_addr(mem_0_15_R0_addr),
    .R0_clk(mem_0_15_R0_clk),
    .R0_data(mem_0_15_R0_data),
    .R0_en(mem_0_15_R0_en)
  );
  split_mem_0_ext mem_0_16 (
    .W0_addr(mem_0_16_W0_addr),
    .W0_clk(mem_0_16_W0_clk),
    .W0_data(mem_0_16_W0_data),
    .W0_en(mem_0_16_W0_en),
    .W0_mask(mem_0_16_W0_mask),
    .R0_addr(mem_0_16_R0_addr),
    .R0_clk(mem_0_16_R0_clk),
    .R0_data(mem_0_16_R0_data),
    .R0_en(mem_0_16_R0_en)
  );
  split_mem_0_ext mem_0_17 (
    .W0_addr(mem_0_17_W0_addr),
    .W0_clk(mem_0_17_W0_clk),
    .W0_data(mem_0_17_W0_data),
    .W0_en(mem_0_17_W0_en),
    .W0_mask(mem_0_17_W0_mask),
    .R0_addr(mem_0_17_R0_addr),
    .R0_clk(mem_0_17_R0_clk),
    .R0_data(mem_0_17_R0_data),
    .R0_en(mem_0_17_R0_en)
  );
  split_mem_0_ext mem_0_18 (
    .W0_addr(mem_0_18_W0_addr),
    .W0_clk(mem_0_18_W0_clk),
    .W0_data(mem_0_18_W0_data),
    .W0_en(mem_0_18_W0_en),
    .W0_mask(mem_0_18_W0_mask),
    .R0_addr(mem_0_18_R0_addr),
    .R0_clk(mem_0_18_R0_clk),
    .R0_data(mem_0_18_R0_data),
    .R0_en(mem_0_18_R0_en)
  );
  split_mem_0_ext mem_0_19 (
    .W0_addr(mem_0_19_W0_addr),
    .W0_clk(mem_0_19_W0_clk),
    .W0_data(mem_0_19_W0_data),
    .W0_en(mem_0_19_W0_en),
    .W0_mask(mem_0_19_W0_mask),
    .R0_addr(mem_0_19_R0_addr),
    .R0_clk(mem_0_19_R0_clk),
    .R0_data(mem_0_19_R0_data),
    .R0_en(mem_0_19_R0_en)
  );
  split_mem_0_ext mem_0_20 (
    .W0_addr(mem_0_20_W0_addr),
    .W0_clk(mem_0_20_W0_clk),
    .W0_data(mem_0_20_W0_data),
    .W0_en(mem_0_20_W0_en),
    .W0_mask(mem_0_20_W0_mask),
    .R0_addr(mem_0_20_R0_addr),
    .R0_clk(mem_0_20_R0_clk),
    .R0_data(mem_0_20_R0_data),
    .R0_en(mem_0_20_R0_en)
  );
  split_mem_0_ext mem_0_21 (
    .W0_addr(mem_0_21_W0_addr),
    .W0_clk(mem_0_21_W0_clk),
    .W0_data(mem_0_21_W0_data),
    .W0_en(mem_0_21_W0_en),
    .W0_mask(mem_0_21_W0_mask),
    .R0_addr(mem_0_21_R0_addr),
    .R0_clk(mem_0_21_R0_clk),
    .R0_data(mem_0_21_R0_data),
    .R0_en(mem_0_21_R0_en)
  );
  split_mem_0_ext mem_0_22 (
    .W0_addr(mem_0_22_W0_addr),
    .W0_clk(mem_0_22_W0_clk),
    .W0_data(mem_0_22_W0_data),
    .W0_en(mem_0_22_W0_en),
    .W0_mask(mem_0_22_W0_mask),
    .R0_addr(mem_0_22_R0_addr),
    .R0_clk(mem_0_22_R0_clk),
    .R0_data(mem_0_22_R0_data),
    .R0_en(mem_0_22_R0_en)
  );
  split_mem_0_ext mem_0_23 (
    .W0_addr(mem_0_23_W0_addr),
    .W0_clk(mem_0_23_W0_clk),
    .W0_data(mem_0_23_W0_data),
    .W0_en(mem_0_23_W0_en),
    .W0_mask(mem_0_23_W0_mask),
    .R0_addr(mem_0_23_R0_addr),
    .R0_clk(mem_0_23_R0_clk),
    .R0_data(mem_0_23_R0_data),
    .R0_en(mem_0_23_R0_en)
  );
  split_mem_0_ext mem_0_24 (
    .W0_addr(mem_0_24_W0_addr),
    .W0_clk(mem_0_24_W0_clk),
    .W0_data(mem_0_24_W0_data),
    .W0_en(mem_0_24_W0_en),
    .W0_mask(mem_0_24_W0_mask),
    .R0_addr(mem_0_24_R0_addr),
    .R0_clk(mem_0_24_R0_clk),
    .R0_data(mem_0_24_R0_data),
    .R0_en(mem_0_24_R0_en)
  );
  split_mem_0_ext mem_0_25 (
    .W0_addr(mem_0_25_W0_addr),
    .W0_clk(mem_0_25_W0_clk),
    .W0_data(mem_0_25_W0_data),
    .W0_en(mem_0_25_W0_en),
    .W0_mask(mem_0_25_W0_mask),
    .R0_addr(mem_0_25_R0_addr),
    .R0_clk(mem_0_25_R0_clk),
    .R0_data(mem_0_25_R0_data),
    .R0_en(mem_0_25_R0_en)
  );
  split_mem_0_ext mem_0_26 (
    .W0_addr(mem_0_26_W0_addr),
    .W0_clk(mem_0_26_W0_clk),
    .W0_data(mem_0_26_W0_data),
    .W0_en(mem_0_26_W0_en),
    .W0_mask(mem_0_26_W0_mask),
    .R0_addr(mem_0_26_R0_addr),
    .R0_clk(mem_0_26_R0_clk),
    .R0_data(mem_0_26_R0_data),
    .R0_en(mem_0_26_R0_en)
  );
  split_mem_0_ext mem_0_27 (
    .W0_addr(mem_0_27_W0_addr),
    .W0_clk(mem_0_27_W0_clk),
    .W0_data(mem_0_27_W0_data),
    .W0_en(mem_0_27_W0_en),
    .W0_mask(mem_0_27_W0_mask),
    .R0_addr(mem_0_27_R0_addr),
    .R0_clk(mem_0_27_R0_clk),
    .R0_data(mem_0_27_R0_data),
    .R0_en(mem_0_27_R0_en)
  );
  split_mem_0_ext mem_0_28 (
    .W0_addr(mem_0_28_W0_addr),
    .W0_clk(mem_0_28_W0_clk),
    .W0_data(mem_0_28_W0_data),
    .W0_en(mem_0_28_W0_en),
    .W0_mask(mem_0_28_W0_mask),
    .R0_addr(mem_0_28_R0_addr),
    .R0_clk(mem_0_28_R0_clk),
    .R0_data(mem_0_28_R0_data),
    .R0_en(mem_0_28_R0_en)
  );
  split_mem_0_ext mem_0_29 (
    .W0_addr(mem_0_29_W0_addr),
    .W0_clk(mem_0_29_W0_clk),
    .W0_data(mem_0_29_W0_data),
    .W0_en(mem_0_29_W0_en),
    .W0_mask(mem_0_29_W0_mask),
    .R0_addr(mem_0_29_R0_addr),
    .R0_clk(mem_0_29_R0_clk),
    .R0_data(mem_0_29_R0_data),
    .R0_en(mem_0_29_R0_en)
  );
  split_mem_0_ext mem_0_30 (
    .W0_addr(mem_0_30_W0_addr),
    .W0_clk(mem_0_30_W0_clk),
    .W0_data(mem_0_30_W0_data),
    .W0_en(mem_0_30_W0_en),
    .W0_mask(mem_0_30_W0_mask),
    .R0_addr(mem_0_30_R0_addr),
    .R0_clk(mem_0_30_R0_clk),
    .R0_data(mem_0_30_R0_data),
    .R0_en(mem_0_30_R0_en)
  );
  split_mem_0_ext mem_0_31 (
    .W0_addr(mem_0_31_W0_addr),
    .W0_clk(mem_0_31_W0_clk),
    .W0_data(mem_0_31_W0_data),
    .W0_en(mem_0_31_W0_en),
    .W0_mask(mem_0_31_W0_mask),
    .R0_addr(mem_0_31_R0_addr),
    .R0_clk(mem_0_31_R0_clk),
    .R0_data(mem_0_31_R0_data),
    .R0_en(mem_0_31_R0_en)
  );
  split_mem_0_ext mem_0_32 (
    .W0_addr(mem_0_32_W0_addr),
    .W0_clk(mem_0_32_W0_clk),
    .W0_data(mem_0_32_W0_data),
    .W0_en(mem_0_32_W0_en),
    .W0_mask(mem_0_32_W0_mask),
    .R0_addr(mem_0_32_R0_addr),
    .R0_clk(mem_0_32_R0_clk),
    .R0_data(mem_0_32_R0_data),
    .R0_en(mem_0_32_R0_en)
  );
  split_mem_0_ext mem_0_33 (
    .W0_addr(mem_0_33_W0_addr),
    .W0_clk(mem_0_33_W0_clk),
    .W0_data(mem_0_33_W0_data),
    .W0_en(mem_0_33_W0_en),
    .W0_mask(mem_0_33_W0_mask),
    .R0_addr(mem_0_33_R0_addr),
    .R0_clk(mem_0_33_R0_clk),
    .R0_data(mem_0_33_R0_data),
    .R0_en(mem_0_33_R0_en)
  );
  split_mem_0_ext mem_0_34 (
    .W0_addr(mem_0_34_W0_addr),
    .W0_clk(mem_0_34_W0_clk),
    .W0_data(mem_0_34_W0_data),
    .W0_en(mem_0_34_W0_en),
    .W0_mask(mem_0_34_W0_mask),
    .R0_addr(mem_0_34_R0_addr),
    .R0_clk(mem_0_34_R0_clk),
    .R0_data(mem_0_34_R0_data),
    .R0_en(mem_0_34_R0_en)
  );
  split_mem_0_ext mem_0_35 (
    .W0_addr(mem_0_35_W0_addr),
    .W0_clk(mem_0_35_W0_clk),
    .W0_data(mem_0_35_W0_data),
    .W0_en(mem_0_35_W0_en),
    .W0_mask(mem_0_35_W0_mask),
    .R0_addr(mem_0_35_R0_addr),
    .R0_clk(mem_0_35_R0_clk),
    .R0_data(mem_0_35_R0_data),
    .R0_en(mem_0_35_R0_en)
  );
  split_mem_0_ext mem_0_36 (
    .W0_addr(mem_0_36_W0_addr),
    .W0_clk(mem_0_36_W0_clk),
    .W0_data(mem_0_36_W0_data),
    .W0_en(mem_0_36_W0_en),
    .W0_mask(mem_0_36_W0_mask),
    .R0_addr(mem_0_36_R0_addr),
    .R0_clk(mem_0_36_R0_clk),
    .R0_data(mem_0_36_R0_data),
    .R0_en(mem_0_36_R0_en)
  );
  split_mem_0_ext mem_0_37 (
    .W0_addr(mem_0_37_W0_addr),
    .W0_clk(mem_0_37_W0_clk),
    .W0_data(mem_0_37_W0_data),
    .W0_en(mem_0_37_W0_en),
    .W0_mask(mem_0_37_W0_mask),
    .R0_addr(mem_0_37_R0_addr),
    .R0_clk(mem_0_37_R0_clk),
    .R0_data(mem_0_37_R0_data),
    .R0_en(mem_0_37_R0_en)
  );
  split_mem_0_ext mem_0_38 (
    .W0_addr(mem_0_38_W0_addr),
    .W0_clk(mem_0_38_W0_clk),
    .W0_data(mem_0_38_W0_data),
    .W0_en(mem_0_38_W0_en),
    .W0_mask(mem_0_38_W0_mask),
    .R0_addr(mem_0_38_R0_addr),
    .R0_clk(mem_0_38_R0_clk),
    .R0_data(mem_0_38_R0_data),
    .R0_en(mem_0_38_R0_en)
  );
  split_mem_0_ext mem_0_39 (
    .W0_addr(mem_0_39_W0_addr),
    .W0_clk(mem_0_39_W0_clk),
    .W0_data(mem_0_39_W0_data),
    .W0_en(mem_0_39_W0_en),
    .W0_mask(mem_0_39_W0_mask),
    .R0_addr(mem_0_39_R0_addr),
    .R0_clk(mem_0_39_R0_clk),
    .R0_data(mem_0_39_R0_data),
    .R0_en(mem_0_39_R0_en)
  );
  split_mem_0_ext mem_0_40 (
    .W0_addr(mem_0_40_W0_addr),
    .W0_clk(mem_0_40_W0_clk),
    .W0_data(mem_0_40_W0_data),
    .W0_en(mem_0_40_W0_en),
    .W0_mask(mem_0_40_W0_mask),
    .R0_addr(mem_0_40_R0_addr),
    .R0_clk(mem_0_40_R0_clk),
    .R0_data(mem_0_40_R0_data),
    .R0_en(mem_0_40_R0_en)
  );
  split_mem_0_ext mem_0_41 (
    .W0_addr(mem_0_41_W0_addr),
    .W0_clk(mem_0_41_W0_clk),
    .W0_data(mem_0_41_W0_data),
    .W0_en(mem_0_41_W0_en),
    .W0_mask(mem_0_41_W0_mask),
    .R0_addr(mem_0_41_R0_addr),
    .R0_clk(mem_0_41_R0_clk),
    .R0_data(mem_0_41_R0_data),
    .R0_en(mem_0_41_R0_en)
  );
  split_mem_0_ext mem_0_42 (
    .W0_addr(mem_0_42_W0_addr),
    .W0_clk(mem_0_42_W0_clk),
    .W0_data(mem_0_42_W0_data),
    .W0_en(mem_0_42_W0_en),
    .W0_mask(mem_0_42_W0_mask),
    .R0_addr(mem_0_42_R0_addr),
    .R0_clk(mem_0_42_R0_clk),
    .R0_data(mem_0_42_R0_data),
    .R0_en(mem_0_42_R0_en)
  );
  split_mem_0_ext mem_0_43 (
    .W0_addr(mem_0_43_W0_addr),
    .W0_clk(mem_0_43_W0_clk),
    .W0_data(mem_0_43_W0_data),
    .W0_en(mem_0_43_W0_en),
    .W0_mask(mem_0_43_W0_mask),
    .R0_addr(mem_0_43_R0_addr),
    .R0_clk(mem_0_43_R0_clk),
    .R0_data(mem_0_43_R0_data),
    .R0_en(mem_0_43_R0_en)
  );
  split_mem_0_ext mem_0_44 (
    .W0_addr(mem_0_44_W0_addr),
    .W0_clk(mem_0_44_W0_clk),
    .W0_data(mem_0_44_W0_data),
    .W0_en(mem_0_44_W0_en),
    .W0_mask(mem_0_44_W0_mask),
    .R0_addr(mem_0_44_R0_addr),
    .R0_clk(mem_0_44_R0_clk),
    .R0_data(mem_0_44_R0_data),
    .R0_en(mem_0_44_R0_en)
  );
  split_mem_0_ext mem_0_45 (
    .W0_addr(mem_0_45_W0_addr),
    .W0_clk(mem_0_45_W0_clk),
    .W0_data(mem_0_45_W0_data),
    .W0_en(mem_0_45_W0_en),
    .W0_mask(mem_0_45_W0_mask),
    .R0_addr(mem_0_45_R0_addr),
    .R0_clk(mem_0_45_R0_clk),
    .R0_data(mem_0_45_R0_data),
    .R0_en(mem_0_45_R0_en)
  );
  split_mem_0_ext mem_0_46 (
    .W0_addr(mem_0_46_W0_addr),
    .W0_clk(mem_0_46_W0_clk),
    .W0_data(mem_0_46_W0_data),
    .W0_en(mem_0_46_W0_en),
    .W0_mask(mem_0_46_W0_mask),
    .R0_addr(mem_0_46_R0_addr),
    .R0_clk(mem_0_46_R0_clk),
    .R0_data(mem_0_46_R0_data),
    .R0_en(mem_0_46_R0_en)
  );
  split_mem_0_ext mem_0_47 (
    .W0_addr(mem_0_47_W0_addr),
    .W0_clk(mem_0_47_W0_clk),
    .W0_data(mem_0_47_W0_data),
    .W0_en(mem_0_47_W0_en),
    .W0_mask(mem_0_47_W0_mask),
    .R0_addr(mem_0_47_R0_addr),
    .R0_clk(mem_0_47_R0_clk),
    .R0_data(mem_0_47_R0_data),
    .R0_en(mem_0_47_R0_en)
  );
  split_mem_0_ext mem_0_48 (
    .W0_addr(mem_0_48_W0_addr),
    .W0_clk(mem_0_48_W0_clk),
    .W0_data(mem_0_48_W0_data),
    .W0_en(mem_0_48_W0_en),
    .W0_mask(mem_0_48_W0_mask),
    .R0_addr(mem_0_48_R0_addr),
    .R0_clk(mem_0_48_R0_clk),
    .R0_data(mem_0_48_R0_data),
    .R0_en(mem_0_48_R0_en)
  );
  split_mem_0_ext mem_0_49 (
    .W0_addr(mem_0_49_W0_addr),
    .W0_clk(mem_0_49_W0_clk),
    .W0_data(mem_0_49_W0_data),
    .W0_en(mem_0_49_W0_en),
    .W0_mask(mem_0_49_W0_mask),
    .R0_addr(mem_0_49_R0_addr),
    .R0_clk(mem_0_49_R0_clk),
    .R0_data(mem_0_49_R0_data),
    .R0_en(mem_0_49_R0_en)
  );
  split_mem_0_ext mem_0_50 (
    .W0_addr(mem_0_50_W0_addr),
    .W0_clk(mem_0_50_W0_clk),
    .W0_data(mem_0_50_W0_data),
    .W0_en(mem_0_50_W0_en),
    .W0_mask(mem_0_50_W0_mask),
    .R0_addr(mem_0_50_R0_addr),
    .R0_clk(mem_0_50_R0_clk),
    .R0_data(mem_0_50_R0_data),
    .R0_en(mem_0_50_R0_en)
  );
  split_mem_0_ext mem_0_51 (
    .W0_addr(mem_0_51_W0_addr),
    .W0_clk(mem_0_51_W0_clk),
    .W0_data(mem_0_51_W0_data),
    .W0_en(mem_0_51_W0_en),
    .W0_mask(mem_0_51_W0_mask),
    .R0_addr(mem_0_51_R0_addr),
    .R0_clk(mem_0_51_R0_clk),
    .R0_data(mem_0_51_R0_data),
    .R0_en(mem_0_51_R0_en)
  );
  split_mem_0_ext mem_0_52 (
    .W0_addr(mem_0_52_W0_addr),
    .W0_clk(mem_0_52_W0_clk),
    .W0_data(mem_0_52_W0_data),
    .W0_en(mem_0_52_W0_en),
    .W0_mask(mem_0_52_W0_mask),
    .R0_addr(mem_0_52_R0_addr),
    .R0_clk(mem_0_52_R0_clk),
    .R0_data(mem_0_52_R0_data),
    .R0_en(mem_0_52_R0_en)
  );
  split_mem_0_ext mem_0_53 (
    .W0_addr(mem_0_53_W0_addr),
    .W0_clk(mem_0_53_W0_clk),
    .W0_data(mem_0_53_W0_data),
    .W0_en(mem_0_53_W0_en),
    .W0_mask(mem_0_53_W0_mask),
    .R0_addr(mem_0_53_R0_addr),
    .R0_clk(mem_0_53_R0_clk),
    .R0_data(mem_0_53_R0_data),
    .R0_en(mem_0_53_R0_en)
  );
  split_mem_0_ext mem_0_54 (
    .W0_addr(mem_0_54_W0_addr),
    .W0_clk(mem_0_54_W0_clk),
    .W0_data(mem_0_54_W0_data),
    .W0_en(mem_0_54_W0_en),
    .W0_mask(mem_0_54_W0_mask),
    .R0_addr(mem_0_54_R0_addr),
    .R0_clk(mem_0_54_R0_clk),
    .R0_data(mem_0_54_R0_data),
    .R0_en(mem_0_54_R0_en)
  );
  split_mem_0_ext mem_0_55 (
    .W0_addr(mem_0_55_W0_addr),
    .W0_clk(mem_0_55_W0_clk),
    .W0_data(mem_0_55_W0_data),
    .W0_en(mem_0_55_W0_en),
    .W0_mask(mem_0_55_W0_mask),
    .R0_addr(mem_0_55_R0_addr),
    .R0_clk(mem_0_55_R0_clk),
    .R0_data(mem_0_55_R0_data),
    .R0_en(mem_0_55_R0_en)
  );
  split_mem_0_ext mem_0_56 (
    .W0_addr(mem_0_56_W0_addr),
    .W0_clk(mem_0_56_W0_clk),
    .W0_data(mem_0_56_W0_data),
    .W0_en(mem_0_56_W0_en),
    .W0_mask(mem_0_56_W0_mask),
    .R0_addr(mem_0_56_R0_addr),
    .R0_clk(mem_0_56_R0_clk),
    .R0_data(mem_0_56_R0_data),
    .R0_en(mem_0_56_R0_en)
  );
  split_mem_0_ext mem_0_57 (
    .W0_addr(mem_0_57_W0_addr),
    .W0_clk(mem_0_57_W0_clk),
    .W0_data(mem_0_57_W0_data),
    .W0_en(mem_0_57_W0_en),
    .W0_mask(mem_0_57_W0_mask),
    .R0_addr(mem_0_57_R0_addr),
    .R0_clk(mem_0_57_R0_clk),
    .R0_data(mem_0_57_R0_data),
    .R0_en(mem_0_57_R0_en)
  );
  split_mem_0_ext mem_0_58 (
    .W0_addr(mem_0_58_W0_addr),
    .W0_clk(mem_0_58_W0_clk),
    .W0_data(mem_0_58_W0_data),
    .W0_en(mem_0_58_W0_en),
    .W0_mask(mem_0_58_W0_mask),
    .R0_addr(mem_0_58_R0_addr),
    .R0_clk(mem_0_58_R0_clk),
    .R0_data(mem_0_58_R0_data),
    .R0_en(mem_0_58_R0_en)
  );
  split_mem_0_ext mem_0_59 (
    .W0_addr(mem_0_59_W0_addr),
    .W0_clk(mem_0_59_W0_clk),
    .W0_data(mem_0_59_W0_data),
    .W0_en(mem_0_59_W0_en),
    .W0_mask(mem_0_59_W0_mask),
    .R0_addr(mem_0_59_R0_addr),
    .R0_clk(mem_0_59_R0_clk),
    .R0_data(mem_0_59_R0_data),
    .R0_en(mem_0_59_R0_en)
  );
  split_mem_0_ext mem_0_60 (
    .W0_addr(mem_0_60_W0_addr),
    .W0_clk(mem_0_60_W0_clk),
    .W0_data(mem_0_60_W0_data),
    .W0_en(mem_0_60_W0_en),
    .W0_mask(mem_0_60_W0_mask),
    .R0_addr(mem_0_60_R0_addr),
    .R0_clk(mem_0_60_R0_clk),
    .R0_data(mem_0_60_R0_data),
    .R0_en(mem_0_60_R0_en)
  );
  split_mem_0_ext mem_0_61 (
    .W0_addr(mem_0_61_W0_addr),
    .W0_clk(mem_0_61_W0_clk),
    .W0_data(mem_0_61_W0_data),
    .W0_en(mem_0_61_W0_en),
    .W0_mask(mem_0_61_W0_mask),
    .R0_addr(mem_0_61_R0_addr),
    .R0_clk(mem_0_61_R0_clk),
    .R0_data(mem_0_61_R0_data),
    .R0_en(mem_0_61_R0_en)
  );
  split_mem_0_ext mem_0_62 (
    .W0_addr(mem_0_62_W0_addr),
    .W0_clk(mem_0_62_W0_clk),
    .W0_data(mem_0_62_W0_data),
    .W0_en(mem_0_62_W0_en),
    .W0_mask(mem_0_62_W0_mask),
    .R0_addr(mem_0_62_R0_addr),
    .R0_clk(mem_0_62_R0_clk),
    .R0_data(mem_0_62_R0_data),
    .R0_en(mem_0_62_R0_en)
  );
  split_mem_0_ext mem_0_63 (
    .W0_addr(mem_0_63_W0_addr),
    .W0_clk(mem_0_63_W0_clk),
    .W0_data(mem_0_63_W0_data),
    .W0_en(mem_0_63_W0_en),
    .W0_mask(mem_0_63_W0_mask),
    .R0_addr(mem_0_63_R0_addr),
    .R0_clk(mem_0_63_R0_clk),
    .R0_data(mem_0_63_R0_data),
    .R0_en(mem_0_63_R0_en)
  );
  split_mem_0_ext mem_0_64 (
    .W0_addr(mem_0_64_W0_addr),
    .W0_clk(mem_0_64_W0_clk),
    .W0_data(mem_0_64_W0_data),
    .W0_en(mem_0_64_W0_en),
    .W0_mask(mem_0_64_W0_mask),
    .R0_addr(mem_0_64_R0_addr),
    .R0_clk(mem_0_64_R0_clk),
    .R0_data(mem_0_64_R0_data),
    .R0_en(mem_0_64_R0_en)
  );
  split_mem_0_ext mem_0_65 (
    .W0_addr(mem_0_65_W0_addr),
    .W0_clk(mem_0_65_W0_clk),
    .W0_data(mem_0_65_W0_data),
    .W0_en(mem_0_65_W0_en),
    .W0_mask(mem_0_65_W0_mask),
    .R0_addr(mem_0_65_R0_addr),
    .R0_clk(mem_0_65_R0_clk),
    .R0_data(mem_0_65_R0_data),
    .R0_en(mem_0_65_R0_en)
  );
  split_mem_0_ext mem_0_66 (
    .W0_addr(mem_0_66_W0_addr),
    .W0_clk(mem_0_66_W0_clk),
    .W0_data(mem_0_66_W0_data),
    .W0_en(mem_0_66_W0_en),
    .W0_mask(mem_0_66_W0_mask),
    .R0_addr(mem_0_66_R0_addr),
    .R0_clk(mem_0_66_R0_clk),
    .R0_data(mem_0_66_R0_data),
    .R0_en(mem_0_66_R0_en)
  );
  split_mem_0_ext mem_0_67 (
    .W0_addr(mem_0_67_W0_addr),
    .W0_clk(mem_0_67_W0_clk),
    .W0_data(mem_0_67_W0_data),
    .W0_en(mem_0_67_W0_en),
    .W0_mask(mem_0_67_W0_mask),
    .R0_addr(mem_0_67_R0_addr),
    .R0_clk(mem_0_67_R0_clk),
    .R0_data(mem_0_67_R0_data),
    .R0_en(mem_0_67_R0_en)
  );
  split_mem_0_ext mem_0_68 (
    .W0_addr(mem_0_68_W0_addr),
    .W0_clk(mem_0_68_W0_clk),
    .W0_data(mem_0_68_W0_data),
    .W0_en(mem_0_68_W0_en),
    .W0_mask(mem_0_68_W0_mask),
    .R0_addr(mem_0_68_R0_addr),
    .R0_clk(mem_0_68_R0_clk),
    .R0_data(mem_0_68_R0_data),
    .R0_en(mem_0_68_R0_en)
  );
  split_mem_0_ext mem_0_69 (
    .W0_addr(mem_0_69_W0_addr),
    .W0_clk(mem_0_69_W0_clk),
    .W0_data(mem_0_69_W0_data),
    .W0_en(mem_0_69_W0_en),
    .W0_mask(mem_0_69_W0_mask),
    .R0_addr(mem_0_69_R0_addr),
    .R0_clk(mem_0_69_R0_clk),
    .R0_data(mem_0_69_R0_data),
    .R0_en(mem_0_69_R0_en)
  );
  split_mem_0_ext mem_0_70 (
    .W0_addr(mem_0_70_W0_addr),
    .W0_clk(mem_0_70_W0_clk),
    .W0_data(mem_0_70_W0_data),
    .W0_en(mem_0_70_W0_en),
    .W0_mask(mem_0_70_W0_mask),
    .R0_addr(mem_0_70_R0_addr),
    .R0_clk(mem_0_70_R0_clk),
    .R0_data(mem_0_70_R0_data),
    .R0_en(mem_0_70_R0_en)
  );
  split_mem_0_ext mem_0_71 (
    .W0_addr(mem_0_71_W0_addr),
    .W0_clk(mem_0_71_W0_clk),
    .W0_data(mem_0_71_W0_data),
    .W0_en(mem_0_71_W0_en),
    .W0_mask(mem_0_71_W0_mask),
    .R0_addr(mem_0_71_R0_addr),
    .R0_clk(mem_0_71_R0_clk),
    .R0_data(mem_0_71_R0_data),
    .R0_en(mem_0_71_R0_en)
  );
  split_mem_0_ext mem_0_72 (
    .W0_addr(mem_0_72_W0_addr),
    .W0_clk(mem_0_72_W0_clk),
    .W0_data(mem_0_72_W0_data),
    .W0_en(mem_0_72_W0_en),
    .W0_mask(mem_0_72_W0_mask),
    .R0_addr(mem_0_72_R0_addr),
    .R0_clk(mem_0_72_R0_clk),
    .R0_data(mem_0_72_R0_data),
    .R0_en(mem_0_72_R0_en)
  );
  split_mem_0_ext mem_0_73 (
    .W0_addr(mem_0_73_W0_addr),
    .W0_clk(mem_0_73_W0_clk),
    .W0_data(mem_0_73_W0_data),
    .W0_en(mem_0_73_W0_en),
    .W0_mask(mem_0_73_W0_mask),
    .R0_addr(mem_0_73_R0_addr),
    .R0_clk(mem_0_73_R0_clk),
    .R0_data(mem_0_73_R0_data),
    .R0_en(mem_0_73_R0_en)
  );
  split_mem_0_ext mem_0_74 (
    .W0_addr(mem_0_74_W0_addr),
    .W0_clk(mem_0_74_W0_clk),
    .W0_data(mem_0_74_W0_data),
    .W0_en(mem_0_74_W0_en),
    .W0_mask(mem_0_74_W0_mask),
    .R0_addr(mem_0_74_R0_addr),
    .R0_clk(mem_0_74_R0_clk),
    .R0_data(mem_0_74_R0_data),
    .R0_en(mem_0_74_R0_en)
  );
  split_mem_0_ext mem_0_75 (
    .W0_addr(mem_0_75_W0_addr),
    .W0_clk(mem_0_75_W0_clk),
    .W0_data(mem_0_75_W0_data),
    .W0_en(mem_0_75_W0_en),
    .W0_mask(mem_0_75_W0_mask),
    .R0_addr(mem_0_75_R0_addr),
    .R0_clk(mem_0_75_R0_clk),
    .R0_data(mem_0_75_R0_data),
    .R0_en(mem_0_75_R0_en)
  );
  split_mem_0_ext mem_0_76 (
    .W0_addr(mem_0_76_W0_addr),
    .W0_clk(mem_0_76_W0_clk),
    .W0_data(mem_0_76_W0_data),
    .W0_en(mem_0_76_W0_en),
    .W0_mask(mem_0_76_W0_mask),
    .R0_addr(mem_0_76_R0_addr),
    .R0_clk(mem_0_76_R0_clk),
    .R0_data(mem_0_76_R0_data),
    .R0_en(mem_0_76_R0_en)
  );
  split_mem_0_ext mem_0_77 (
    .W0_addr(mem_0_77_W0_addr),
    .W0_clk(mem_0_77_W0_clk),
    .W0_data(mem_0_77_W0_data),
    .W0_en(mem_0_77_W0_en),
    .W0_mask(mem_0_77_W0_mask),
    .R0_addr(mem_0_77_R0_addr),
    .R0_clk(mem_0_77_R0_clk),
    .R0_data(mem_0_77_R0_data),
    .R0_en(mem_0_77_R0_en)
  );
  split_mem_0_ext mem_0_78 (
    .W0_addr(mem_0_78_W0_addr),
    .W0_clk(mem_0_78_W0_clk),
    .W0_data(mem_0_78_W0_data),
    .W0_en(mem_0_78_W0_en),
    .W0_mask(mem_0_78_W0_mask),
    .R0_addr(mem_0_78_R0_addr),
    .R0_clk(mem_0_78_R0_clk),
    .R0_data(mem_0_78_R0_data),
    .R0_en(mem_0_78_R0_en)
  );
  split_mem_0_ext mem_0_79 (
    .W0_addr(mem_0_79_W0_addr),
    .W0_clk(mem_0_79_W0_clk),
    .W0_data(mem_0_79_W0_data),
    .W0_en(mem_0_79_W0_en),
    .W0_mask(mem_0_79_W0_mask),
    .R0_addr(mem_0_79_R0_addr),
    .R0_clk(mem_0_79_R0_clk),
    .R0_data(mem_0_79_R0_data),
    .R0_en(mem_0_79_R0_en)
  );
  split_mem_0_ext mem_0_80 (
    .W0_addr(mem_0_80_W0_addr),
    .W0_clk(mem_0_80_W0_clk),
    .W0_data(mem_0_80_W0_data),
    .W0_en(mem_0_80_W0_en),
    .W0_mask(mem_0_80_W0_mask),
    .R0_addr(mem_0_80_R0_addr),
    .R0_clk(mem_0_80_R0_clk),
    .R0_data(mem_0_80_R0_data),
    .R0_en(mem_0_80_R0_en)
  );
  split_mem_0_ext mem_0_81 (
    .W0_addr(mem_0_81_W0_addr),
    .W0_clk(mem_0_81_W0_clk),
    .W0_data(mem_0_81_W0_data),
    .W0_en(mem_0_81_W0_en),
    .W0_mask(mem_0_81_W0_mask),
    .R0_addr(mem_0_81_R0_addr),
    .R0_clk(mem_0_81_R0_clk),
    .R0_data(mem_0_81_R0_data),
    .R0_en(mem_0_81_R0_en)
  );
  split_mem_0_ext mem_0_82 (
    .W0_addr(mem_0_82_W0_addr),
    .W0_clk(mem_0_82_W0_clk),
    .W0_data(mem_0_82_W0_data),
    .W0_en(mem_0_82_W0_en),
    .W0_mask(mem_0_82_W0_mask),
    .R0_addr(mem_0_82_R0_addr),
    .R0_clk(mem_0_82_R0_clk),
    .R0_data(mem_0_82_R0_data),
    .R0_en(mem_0_82_R0_en)
  );
  split_mem_0_ext mem_0_83 (
    .W0_addr(mem_0_83_W0_addr),
    .W0_clk(mem_0_83_W0_clk),
    .W0_data(mem_0_83_W0_data),
    .W0_en(mem_0_83_W0_en),
    .W0_mask(mem_0_83_W0_mask),
    .R0_addr(mem_0_83_R0_addr),
    .R0_clk(mem_0_83_R0_clk),
    .R0_data(mem_0_83_R0_data),
    .R0_en(mem_0_83_R0_en)
  );
  split_mem_0_ext mem_0_84 (
    .W0_addr(mem_0_84_W0_addr),
    .W0_clk(mem_0_84_W0_clk),
    .W0_data(mem_0_84_W0_data),
    .W0_en(mem_0_84_W0_en),
    .W0_mask(mem_0_84_W0_mask),
    .R0_addr(mem_0_84_R0_addr),
    .R0_clk(mem_0_84_R0_clk),
    .R0_data(mem_0_84_R0_data),
    .R0_en(mem_0_84_R0_en)
  );
  split_mem_0_ext mem_0_85 (
    .W0_addr(mem_0_85_W0_addr),
    .W0_clk(mem_0_85_W0_clk),
    .W0_data(mem_0_85_W0_data),
    .W0_en(mem_0_85_W0_en),
    .W0_mask(mem_0_85_W0_mask),
    .R0_addr(mem_0_85_R0_addr),
    .R0_clk(mem_0_85_R0_clk),
    .R0_data(mem_0_85_R0_data),
    .R0_en(mem_0_85_R0_en)
  );
  split_mem_0_ext mem_0_86 (
    .W0_addr(mem_0_86_W0_addr),
    .W0_clk(mem_0_86_W0_clk),
    .W0_data(mem_0_86_W0_data),
    .W0_en(mem_0_86_W0_en),
    .W0_mask(mem_0_86_W0_mask),
    .R0_addr(mem_0_86_R0_addr),
    .R0_clk(mem_0_86_R0_clk),
    .R0_data(mem_0_86_R0_data),
    .R0_en(mem_0_86_R0_en)
  );
  split_mem_0_ext mem_0_87 (
    .W0_addr(mem_0_87_W0_addr),
    .W0_clk(mem_0_87_W0_clk),
    .W0_data(mem_0_87_W0_data),
    .W0_en(mem_0_87_W0_en),
    .W0_mask(mem_0_87_W0_mask),
    .R0_addr(mem_0_87_R0_addr),
    .R0_clk(mem_0_87_R0_clk),
    .R0_data(mem_0_87_R0_data),
    .R0_en(mem_0_87_R0_en)
  );
  split_mem_0_ext mem_0_88 (
    .W0_addr(mem_0_88_W0_addr),
    .W0_clk(mem_0_88_W0_clk),
    .W0_data(mem_0_88_W0_data),
    .W0_en(mem_0_88_W0_en),
    .W0_mask(mem_0_88_W0_mask),
    .R0_addr(mem_0_88_R0_addr),
    .R0_clk(mem_0_88_R0_clk),
    .R0_data(mem_0_88_R0_data),
    .R0_en(mem_0_88_R0_en)
  );
  split_mem_0_ext mem_0_89 (
    .W0_addr(mem_0_89_W0_addr),
    .W0_clk(mem_0_89_W0_clk),
    .W0_data(mem_0_89_W0_data),
    .W0_en(mem_0_89_W0_en),
    .W0_mask(mem_0_89_W0_mask),
    .R0_addr(mem_0_89_R0_addr),
    .R0_clk(mem_0_89_R0_clk),
    .R0_data(mem_0_89_R0_data),
    .R0_en(mem_0_89_R0_en)
  );
  split_mem_0_ext mem_0_90 (
    .W0_addr(mem_0_90_W0_addr),
    .W0_clk(mem_0_90_W0_clk),
    .W0_data(mem_0_90_W0_data),
    .W0_en(mem_0_90_W0_en),
    .W0_mask(mem_0_90_W0_mask),
    .R0_addr(mem_0_90_R0_addr),
    .R0_clk(mem_0_90_R0_clk),
    .R0_data(mem_0_90_R0_data),
    .R0_en(mem_0_90_R0_en)
  );
  split_mem_0_ext mem_0_91 (
    .W0_addr(mem_0_91_W0_addr),
    .W0_clk(mem_0_91_W0_clk),
    .W0_data(mem_0_91_W0_data),
    .W0_en(mem_0_91_W0_en),
    .W0_mask(mem_0_91_W0_mask),
    .R0_addr(mem_0_91_R0_addr),
    .R0_clk(mem_0_91_R0_clk),
    .R0_data(mem_0_91_R0_data),
    .R0_en(mem_0_91_R0_en)
  );
  split_mem_0_ext mem_0_92 (
    .W0_addr(mem_0_92_W0_addr),
    .W0_clk(mem_0_92_W0_clk),
    .W0_data(mem_0_92_W0_data),
    .W0_en(mem_0_92_W0_en),
    .W0_mask(mem_0_92_W0_mask),
    .R0_addr(mem_0_92_R0_addr),
    .R0_clk(mem_0_92_R0_clk),
    .R0_data(mem_0_92_R0_data),
    .R0_en(mem_0_92_R0_en)
  );
  split_mem_0_ext mem_0_93 (
    .W0_addr(mem_0_93_W0_addr),
    .W0_clk(mem_0_93_W0_clk),
    .W0_data(mem_0_93_W0_data),
    .W0_en(mem_0_93_W0_en),
    .W0_mask(mem_0_93_W0_mask),
    .R0_addr(mem_0_93_R0_addr),
    .R0_clk(mem_0_93_R0_clk),
    .R0_data(mem_0_93_R0_data),
    .R0_en(mem_0_93_R0_en)
  );
  split_mem_0_ext mem_0_94 (
    .W0_addr(mem_0_94_W0_addr),
    .W0_clk(mem_0_94_W0_clk),
    .W0_data(mem_0_94_W0_data),
    .W0_en(mem_0_94_W0_en),
    .W0_mask(mem_0_94_W0_mask),
    .R0_addr(mem_0_94_R0_addr),
    .R0_clk(mem_0_94_R0_clk),
    .R0_data(mem_0_94_R0_data),
    .R0_en(mem_0_94_R0_en)
  );
  split_mem_0_ext mem_0_95 (
    .W0_addr(mem_0_95_W0_addr),
    .W0_clk(mem_0_95_W0_clk),
    .W0_data(mem_0_95_W0_data),
    .W0_en(mem_0_95_W0_en),
    .W0_mask(mem_0_95_W0_mask),
    .R0_addr(mem_0_95_R0_addr),
    .R0_clk(mem_0_95_R0_clk),
    .R0_data(mem_0_95_R0_data),
    .R0_en(mem_0_95_R0_en)
  );
  split_mem_0_ext mem_0_96 (
    .W0_addr(mem_0_96_W0_addr),
    .W0_clk(mem_0_96_W0_clk),
    .W0_data(mem_0_96_W0_data),
    .W0_en(mem_0_96_W0_en),
    .W0_mask(mem_0_96_W0_mask),
    .R0_addr(mem_0_96_R0_addr),
    .R0_clk(mem_0_96_R0_clk),
    .R0_data(mem_0_96_R0_data),
    .R0_en(mem_0_96_R0_en)
  );
  split_mem_0_ext mem_0_97 (
    .W0_addr(mem_0_97_W0_addr),
    .W0_clk(mem_0_97_W0_clk),
    .W0_data(mem_0_97_W0_data),
    .W0_en(mem_0_97_W0_en),
    .W0_mask(mem_0_97_W0_mask),
    .R0_addr(mem_0_97_R0_addr),
    .R0_clk(mem_0_97_R0_clk),
    .R0_data(mem_0_97_R0_data),
    .R0_en(mem_0_97_R0_en)
  );
  split_mem_0_ext mem_0_98 (
    .W0_addr(mem_0_98_W0_addr),
    .W0_clk(mem_0_98_W0_clk),
    .W0_data(mem_0_98_W0_data),
    .W0_en(mem_0_98_W0_en),
    .W0_mask(mem_0_98_W0_mask),
    .R0_addr(mem_0_98_R0_addr),
    .R0_clk(mem_0_98_R0_clk),
    .R0_data(mem_0_98_R0_data),
    .R0_en(mem_0_98_R0_en)
  );
  split_mem_0_ext mem_0_99 (
    .W0_addr(mem_0_99_W0_addr),
    .W0_clk(mem_0_99_W0_clk),
    .W0_data(mem_0_99_W0_data),
    .W0_en(mem_0_99_W0_en),
    .W0_mask(mem_0_99_W0_mask),
    .R0_addr(mem_0_99_R0_addr),
    .R0_clk(mem_0_99_R0_clk),
    .R0_data(mem_0_99_R0_data),
    .R0_en(mem_0_99_R0_en)
  );
  split_mem_0_ext mem_0_100 (
    .W0_addr(mem_0_100_W0_addr),
    .W0_clk(mem_0_100_W0_clk),
    .W0_data(mem_0_100_W0_data),
    .W0_en(mem_0_100_W0_en),
    .W0_mask(mem_0_100_W0_mask),
    .R0_addr(mem_0_100_R0_addr),
    .R0_clk(mem_0_100_R0_clk),
    .R0_data(mem_0_100_R0_data),
    .R0_en(mem_0_100_R0_en)
  );
  split_mem_0_ext mem_0_101 (
    .W0_addr(mem_0_101_W0_addr),
    .W0_clk(mem_0_101_W0_clk),
    .W0_data(mem_0_101_W0_data),
    .W0_en(mem_0_101_W0_en),
    .W0_mask(mem_0_101_W0_mask),
    .R0_addr(mem_0_101_R0_addr),
    .R0_clk(mem_0_101_R0_clk),
    .R0_data(mem_0_101_R0_data),
    .R0_en(mem_0_101_R0_en)
  );
  split_mem_0_ext mem_0_102 (
    .W0_addr(mem_0_102_W0_addr),
    .W0_clk(mem_0_102_W0_clk),
    .W0_data(mem_0_102_W0_data),
    .W0_en(mem_0_102_W0_en),
    .W0_mask(mem_0_102_W0_mask),
    .R0_addr(mem_0_102_R0_addr),
    .R0_clk(mem_0_102_R0_clk),
    .R0_data(mem_0_102_R0_data),
    .R0_en(mem_0_102_R0_en)
  );
  split_mem_0_ext mem_0_103 (
    .W0_addr(mem_0_103_W0_addr),
    .W0_clk(mem_0_103_W0_clk),
    .W0_data(mem_0_103_W0_data),
    .W0_en(mem_0_103_W0_en),
    .W0_mask(mem_0_103_W0_mask),
    .R0_addr(mem_0_103_R0_addr),
    .R0_clk(mem_0_103_R0_clk),
    .R0_data(mem_0_103_R0_data),
    .R0_en(mem_0_103_R0_en)
  );
  split_mem_0_ext mem_0_104 (
    .W0_addr(mem_0_104_W0_addr),
    .W0_clk(mem_0_104_W0_clk),
    .W0_data(mem_0_104_W0_data),
    .W0_en(mem_0_104_W0_en),
    .W0_mask(mem_0_104_W0_mask),
    .R0_addr(mem_0_104_R0_addr),
    .R0_clk(mem_0_104_R0_clk),
    .R0_data(mem_0_104_R0_data),
    .R0_en(mem_0_104_R0_en)
  );
  split_mem_0_ext mem_0_105 (
    .W0_addr(mem_0_105_W0_addr),
    .W0_clk(mem_0_105_W0_clk),
    .W0_data(mem_0_105_W0_data),
    .W0_en(mem_0_105_W0_en),
    .W0_mask(mem_0_105_W0_mask),
    .R0_addr(mem_0_105_R0_addr),
    .R0_clk(mem_0_105_R0_clk),
    .R0_data(mem_0_105_R0_data),
    .R0_en(mem_0_105_R0_en)
  );
  split_mem_0_ext mem_0_106 (
    .W0_addr(mem_0_106_W0_addr),
    .W0_clk(mem_0_106_W0_clk),
    .W0_data(mem_0_106_W0_data),
    .W0_en(mem_0_106_W0_en),
    .W0_mask(mem_0_106_W0_mask),
    .R0_addr(mem_0_106_R0_addr),
    .R0_clk(mem_0_106_R0_clk),
    .R0_data(mem_0_106_R0_data),
    .R0_en(mem_0_106_R0_en)
  );
  split_mem_0_ext mem_0_107 (
    .W0_addr(mem_0_107_W0_addr),
    .W0_clk(mem_0_107_W0_clk),
    .W0_data(mem_0_107_W0_data),
    .W0_en(mem_0_107_W0_en),
    .W0_mask(mem_0_107_W0_mask),
    .R0_addr(mem_0_107_R0_addr),
    .R0_clk(mem_0_107_R0_clk),
    .R0_data(mem_0_107_R0_data),
    .R0_en(mem_0_107_R0_en)
  );
  split_mem_0_ext mem_0_108 (
    .W0_addr(mem_0_108_W0_addr),
    .W0_clk(mem_0_108_W0_clk),
    .W0_data(mem_0_108_W0_data),
    .W0_en(mem_0_108_W0_en),
    .W0_mask(mem_0_108_W0_mask),
    .R0_addr(mem_0_108_R0_addr),
    .R0_clk(mem_0_108_R0_clk),
    .R0_data(mem_0_108_R0_data),
    .R0_en(mem_0_108_R0_en)
  );
  split_mem_0_ext mem_0_109 (
    .W0_addr(mem_0_109_W0_addr),
    .W0_clk(mem_0_109_W0_clk),
    .W0_data(mem_0_109_W0_data),
    .W0_en(mem_0_109_W0_en),
    .W0_mask(mem_0_109_W0_mask),
    .R0_addr(mem_0_109_R0_addr),
    .R0_clk(mem_0_109_R0_clk),
    .R0_data(mem_0_109_R0_data),
    .R0_en(mem_0_109_R0_en)
  );
  split_mem_0_ext mem_0_110 (
    .W0_addr(mem_0_110_W0_addr),
    .W0_clk(mem_0_110_W0_clk),
    .W0_data(mem_0_110_W0_data),
    .W0_en(mem_0_110_W0_en),
    .W0_mask(mem_0_110_W0_mask),
    .R0_addr(mem_0_110_R0_addr),
    .R0_clk(mem_0_110_R0_clk),
    .R0_data(mem_0_110_R0_data),
    .R0_en(mem_0_110_R0_en)
  );
  split_mem_0_ext mem_0_111 (
    .W0_addr(mem_0_111_W0_addr),
    .W0_clk(mem_0_111_W0_clk),
    .W0_data(mem_0_111_W0_data),
    .W0_en(mem_0_111_W0_en),
    .W0_mask(mem_0_111_W0_mask),
    .R0_addr(mem_0_111_R0_addr),
    .R0_clk(mem_0_111_R0_clk),
    .R0_data(mem_0_111_R0_data),
    .R0_en(mem_0_111_R0_en)
  );
  split_mem_0_ext mem_0_112 (
    .W0_addr(mem_0_112_W0_addr),
    .W0_clk(mem_0_112_W0_clk),
    .W0_data(mem_0_112_W0_data),
    .W0_en(mem_0_112_W0_en),
    .W0_mask(mem_0_112_W0_mask),
    .R0_addr(mem_0_112_R0_addr),
    .R0_clk(mem_0_112_R0_clk),
    .R0_data(mem_0_112_R0_data),
    .R0_en(mem_0_112_R0_en)
  );
  split_mem_0_ext mem_0_113 (
    .W0_addr(mem_0_113_W0_addr),
    .W0_clk(mem_0_113_W0_clk),
    .W0_data(mem_0_113_W0_data),
    .W0_en(mem_0_113_W0_en),
    .W0_mask(mem_0_113_W0_mask),
    .R0_addr(mem_0_113_R0_addr),
    .R0_clk(mem_0_113_R0_clk),
    .R0_data(mem_0_113_R0_data),
    .R0_en(mem_0_113_R0_en)
  );
  split_mem_0_ext mem_0_114 (
    .W0_addr(mem_0_114_W0_addr),
    .W0_clk(mem_0_114_W0_clk),
    .W0_data(mem_0_114_W0_data),
    .W0_en(mem_0_114_W0_en),
    .W0_mask(mem_0_114_W0_mask),
    .R0_addr(mem_0_114_R0_addr),
    .R0_clk(mem_0_114_R0_clk),
    .R0_data(mem_0_114_R0_data),
    .R0_en(mem_0_114_R0_en)
  );
  split_mem_0_ext mem_0_115 (
    .W0_addr(mem_0_115_W0_addr),
    .W0_clk(mem_0_115_W0_clk),
    .W0_data(mem_0_115_W0_data),
    .W0_en(mem_0_115_W0_en),
    .W0_mask(mem_0_115_W0_mask),
    .R0_addr(mem_0_115_R0_addr),
    .R0_clk(mem_0_115_R0_clk),
    .R0_data(mem_0_115_R0_data),
    .R0_en(mem_0_115_R0_en)
  );
  split_mem_0_ext mem_0_116 (
    .W0_addr(mem_0_116_W0_addr),
    .W0_clk(mem_0_116_W0_clk),
    .W0_data(mem_0_116_W0_data),
    .W0_en(mem_0_116_W0_en),
    .W0_mask(mem_0_116_W0_mask),
    .R0_addr(mem_0_116_R0_addr),
    .R0_clk(mem_0_116_R0_clk),
    .R0_data(mem_0_116_R0_data),
    .R0_en(mem_0_116_R0_en)
  );
  split_mem_0_ext mem_0_117 (
    .W0_addr(mem_0_117_W0_addr),
    .W0_clk(mem_0_117_W0_clk),
    .W0_data(mem_0_117_W0_data),
    .W0_en(mem_0_117_W0_en),
    .W0_mask(mem_0_117_W0_mask),
    .R0_addr(mem_0_117_R0_addr),
    .R0_clk(mem_0_117_R0_clk),
    .R0_data(mem_0_117_R0_data),
    .R0_en(mem_0_117_R0_en)
  );
  split_mem_0_ext mem_0_118 (
    .W0_addr(mem_0_118_W0_addr),
    .W0_clk(mem_0_118_W0_clk),
    .W0_data(mem_0_118_W0_data),
    .W0_en(mem_0_118_W0_en),
    .W0_mask(mem_0_118_W0_mask),
    .R0_addr(mem_0_118_R0_addr),
    .R0_clk(mem_0_118_R0_clk),
    .R0_data(mem_0_118_R0_data),
    .R0_en(mem_0_118_R0_en)
  );
  split_mem_0_ext mem_0_119 (
    .W0_addr(mem_0_119_W0_addr),
    .W0_clk(mem_0_119_W0_clk),
    .W0_data(mem_0_119_W0_data),
    .W0_en(mem_0_119_W0_en),
    .W0_mask(mem_0_119_W0_mask),
    .R0_addr(mem_0_119_R0_addr),
    .R0_clk(mem_0_119_R0_clk),
    .R0_data(mem_0_119_R0_data),
    .R0_en(mem_0_119_R0_en)
  );
  split_mem_0_ext mem_0_120 (
    .W0_addr(mem_0_120_W0_addr),
    .W0_clk(mem_0_120_W0_clk),
    .W0_data(mem_0_120_W0_data),
    .W0_en(mem_0_120_W0_en),
    .W0_mask(mem_0_120_W0_mask),
    .R0_addr(mem_0_120_R0_addr),
    .R0_clk(mem_0_120_R0_clk),
    .R0_data(mem_0_120_R0_data),
    .R0_en(mem_0_120_R0_en)
  );
  split_mem_0_ext mem_0_121 (
    .W0_addr(mem_0_121_W0_addr),
    .W0_clk(mem_0_121_W0_clk),
    .W0_data(mem_0_121_W0_data),
    .W0_en(mem_0_121_W0_en),
    .W0_mask(mem_0_121_W0_mask),
    .R0_addr(mem_0_121_R0_addr),
    .R0_clk(mem_0_121_R0_clk),
    .R0_data(mem_0_121_R0_data),
    .R0_en(mem_0_121_R0_en)
  );
  split_mem_0_ext mem_0_122 (
    .W0_addr(mem_0_122_W0_addr),
    .W0_clk(mem_0_122_W0_clk),
    .W0_data(mem_0_122_W0_data),
    .W0_en(mem_0_122_W0_en),
    .W0_mask(mem_0_122_W0_mask),
    .R0_addr(mem_0_122_R0_addr),
    .R0_clk(mem_0_122_R0_clk),
    .R0_data(mem_0_122_R0_data),
    .R0_en(mem_0_122_R0_en)
  );
  split_mem_0_ext mem_0_123 (
    .W0_addr(mem_0_123_W0_addr),
    .W0_clk(mem_0_123_W0_clk),
    .W0_data(mem_0_123_W0_data),
    .W0_en(mem_0_123_W0_en),
    .W0_mask(mem_0_123_W0_mask),
    .R0_addr(mem_0_123_R0_addr),
    .R0_clk(mem_0_123_R0_clk),
    .R0_data(mem_0_123_R0_data),
    .R0_en(mem_0_123_R0_en)
  );
  split_mem_0_ext mem_0_124 (
    .W0_addr(mem_0_124_W0_addr),
    .W0_clk(mem_0_124_W0_clk),
    .W0_data(mem_0_124_W0_data),
    .W0_en(mem_0_124_W0_en),
    .W0_mask(mem_0_124_W0_mask),
    .R0_addr(mem_0_124_R0_addr),
    .R0_clk(mem_0_124_R0_clk),
    .R0_data(mem_0_124_R0_data),
    .R0_en(mem_0_124_R0_en)
  );
  split_mem_0_ext mem_0_125 (
    .W0_addr(mem_0_125_W0_addr),
    .W0_clk(mem_0_125_W0_clk),
    .W0_data(mem_0_125_W0_data),
    .W0_en(mem_0_125_W0_en),
    .W0_mask(mem_0_125_W0_mask),
    .R0_addr(mem_0_125_R0_addr),
    .R0_clk(mem_0_125_R0_clk),
    .R0_data(mem_0_125_R0_data),
    .R0_en(mem_0_125_R0_en)
  );
  split_mem_0_ext mem_0_126 (
    .W0_addr(mem_0_126_W0_addr),
    .W0_clk(mem_0_126_W0_clk),
    .W0_data(mem_0_126_W0_data),
    .W0_en(mem_0_126_W0_en),
    .W0_mask(mem_0_126_W0_mask),
    .R0_addr(mem_0_126_R0_addr),
    .R0_clk(mem_0_126_R0_clk),
    .R0_data(mem_0_126_R0_data),
    .R0_en(mem_0_126_R0_en)
  );
  split_mem_0_ext mem_0_127 (
    .W0_addr(mem_0_127_W0_addr),
    .W0_clk(mem_0_127_W0_clk),
    .W0_data(mem_0_127_W0_data),
    .W0_en(mem_0_127_W0_en),
    .W0_mask(mem_0_127_W0_mask),
    .R0_addr(mem_0_127_R0_addr),
    .R0_clk(mem_0_127_R0_clk),
    .R0_data(mem_0_127_R0_data),
    .R0_en(mem_0_127_R0_en)
  );
  split_mem_0_ext mem_0_128 (
    .W0_addr(mem_0_128_W0_addr),
    .W0_clk(mem_0_128_W0_clk),
    .W0_data(mem_0_128_W0_data),
    .W0_en(mem_0_128_W0_en),
    .W0_mask(mem_0_128_W0_mask),
    .R0_addr(mem_0_128_R0_addr),
    .R0_clk(mem_0_128_R0_clk),
    .R0_data(mem_0_128_R0_data),
    .R0_en(mem_0_128_R0_en)
  );
  split_mem_0_ext mem_0_129 (
    .W0_addr(mem_0_129_W0_addr),
    .W0_clk(mem_0_129_W0_clk),
    .W0_data(mem_0_129_W0_data),
    .W0_en(mem_0_129_W0_en),
    .W0_mask(mem_0_129_W0_mask),
    .R0_addr(mem_0_129_R0_addr),
    .R0_clk(mem_0_129_R0_clk),
    .R0_data(mem_0_129_R0_data),
    .R0_en(mem_0_129_R0_en)
  );
  split_mem_0_ext mem_0_130 (
    .W0_addr(mem_0_130_W0_addr),
    .W0_clk(mem_0_130_W0_clk),
    .W0_data(mem_0_130_W0_data),
    .W0_en(mem_0_130_W0_en),
    .W0_mask(mem_0_130_W0_mask),
    .R0_addr(mem_0_130_R0_addr),
    .R0_clk(mem_0_130_R0_clk),
    .R0_data(mem_0_130_R0_data),
    .R0_en(mem_0_130_R0_en)
  );
  split_mem_0_ext mem_0_131 (
    .W0_addr(mem_0_131_W0_addr),
    .W0_clk(mem_0_131_W0_clk),
    .W0_data(mem_0_131_W0_data),
    .W0_en(mem_0_131_W0_en),
    .W0_mask(mem_0_131_W0_mask),
    .R0_addr(mem_0_131_R0_addr),
    .R0_clk(mem_0_131_R0_clk),
    .R0_data(mem_0_131_R0_data),
    .R0_en(mem_0_131_R0_en)
  );
  split_mem_0_ext mem_0_132 (
    .W0_addr(mem_0_132_W0_addr),
    .W0_clk(mem_0_132_W0_clk),
    .W0_data(mem_0_132_W0_data),
    .W0_en(mem_0_132_W0_en),
    .W0_mask(mem_0_132_W0_mask),
    .R0_addr(mem_0_132_R0_addr),
    .R0_clk(mem_0_132_R0_clk),
    .R0_data(mem_0_132_R0_data),
    .R0_en(mem_0_132_R0_en)
  );
  split_mem_0_ext mem_0_133 (
    .W0_addr(mem_0_133_W0_addr),
    .W0_clk(mem_0_133_W0_clk),
    .W0_data(mem_0_133_W0_data),
    .W0_en(mem_0_133_W0_en),
    .W0_mask(mem_0_133_W0_mask),
    .R0_addr(mem_0_133_R0_addr),
    .R0_clk(mem_0_133_R0_clk),
    .R0_data(mem_0_133_R0_data),
    .R0_en(mem_0_133_R0_en)
  );
  split_mem_0_ext mem_0_134 (
    .W0_addr(mem_0_134_W0_addr),
    .W0_clk(mem_0_134_W0_clk),
    .W0_data(mem_0_134_W0_data),
    .W0_en(mem_0_134_W0_en),
    .W0_mask(mem_0_134_W0_mask),
    .R0_addr(mem_0_134_R0_addr),
    .R0_clk(mem_0_134_R0_clk),
    .R0_data(mem_0_134_R0_data),
    .R0_en(mem_0_134_R0_en)
  );
  split_mem_0_ext mem_0_135 (
    .W0_addr(mem_0_135_W0_addr),
    .W0_clk(mem_0_135_W0_clk),
    .W0_data(mem_0_135_W0_data),
    .W0_en(mem_0_135_W0_en),
    .W0_mask(mem_0_135_W0_mask),
    .R0_addr(mem_0_135_R0_addr),
    .R0_clk(mem_0_135_R0_clk),
    .R0_data(mem_0_135_R0_data),
    .R0_en(mem_0_135_R0_en)
  );
  split_mem_0_ext mem_0_136 (
    .W0_addr(mem_0_136_W0_addr),
    .W0_clk(mem_0_136_W0_clk),
    .W0_data(mem_0_136_W0_data),
    .W0_en(mem_0_136_W0_en),
    .W0_mask(mem_0_136_W0_mask),
    .R0_addr(mem_0_136_R0_addr),
    .R0_clk(mem_0_136_R0_clk),
    .R0_data(mem_0_136_R0_data),
    .R0_en(mem_0_136_R0_en)
  );
  split_mem_0_ext mem_0_137 (
    .W0_addr(mem_0_137_W0_addr),
    .W0_clk(mem_0_137_W0_clk),
    .W0_data(mem_0_137_W0_data),
    .W0_en(mem_0_137_W0_en),
    .W0_mask(mem_0_137_W0_mask),
    .R0_addr(mem_0_137_R0_addr),
    .R0_clk(mem_0_137_R0_clk),
    .R0_data(mem_0_137_R0_data),
    .R0_en(mem_0_137_R0_en)
  );
  split_mem_0_ext mem_0_138 (
    .W0_addr(mem_0_138_W0_addr),
    .W0_clk(mem_0_138_W0_clk),
    .W0_data(mem_0_138_W0_data),
    .W0_en(mem_0_138_W0_en),
    .W0_mask(mem_0_138_W0_mask),
    .R0_addr(mem_0_138_R0_addr),
    .R0_clk(mem_0_138_R0_clk),
    .R0_data(mem_0_138_R0_data),
    .R0_en(mem_0_138_R0_en)
  );
  split_mem_0_ext mem_0_139 (
    .W0_addr(mem_0_139_W0_addr),
    .W0_clk(mem_0_139_W0_clk),
    .W0_data(mem_0_139_W0_data),
    .W0_en(mem_0_139_W0_en),
    .W0_mask(mem_0_139_W0_mask),
    .R0_addr(mem_0_139_R0_addr),
    .R0_clk(mem_0_139_R0_clk),
    .R0_data(mem_0_139_R0_data),
    .R0_en(mem_0_139_R0_en)
  );
  split_mem_0_ext mem_0_140 (
    .W0_addr(mem_0_140_W0_addr),
    .W0_clk(mem_0_140_W0_clk),
    .W0_data(mem_0_140_W0_data),
    .W0_en(mem_0_140_W0_en),
    .W0_mask(mem_0_140_W0_mask),
    .R0_addr(mem_0_140_R0_addr),
    .R0_clk(mem_0_140_R0_clk),
    .R0_data(mem_0_140_R0_data),
    .R0_en(mem_0_140_R0_en)
  );
  split_mem_0_ext mem_0_141 (
    .W0_addr(mem_0_141_W0_addr),
    .W0_clk(mem_0_141_W0_clk),
    .W0_data(mem_0_141_W0_data),
    .W0_en(mem_0_141_W0_en),
    .W0_mask(mem_0_141_W0_mask),
    .R0_addr(mem_0_141_R0_addr),
    .R0_clk(mem_0_141_R0_clk),
    .R0_data(mem_0_141_R0_data),
    .R0_en(mem_0_141_R0_en)
  );
  split_mem_0_ext mem_0_142 (
    .W0_addr(mem_0_142_W0_addr),
    .W0_clk(mem_0_142_W0_clk),
    .W0_data(mem_0_142_W0_data),
    .W0_en(mem_0_142_W0_en),
    .W0_mask(mem_0_142_W0_mask),
    .R0_addr(mem_0_142_R0_addr),
    .R0_clk(mem_0_142_R0_clk),
    .R0_data(mem_0_142_R0_data),
    .R0_en(mem_0_142_R0_en)
  );
  split_mem_0_ext mem_0_143 (
    .W0_addr(mem_0_143_W0_addr),
    .W0_clk(mem_0_143_W0_clk),
    .W0_data(mem_0_143_W0_data),
    .W0_en(mem_0_143_W0_en),
    .W0_mask(mem_0_143_W0_mask),
    .R0_addr(mem_0_143_R0_addr),
    .R0_clk(mem_0_143_R0_clk),
    .R0_data(mem_0_143_R0_data),
    .R0_en(mem_0_143_R0_en)
  );
  split_mem_0_ext mem_0_144 (
    .W0_addr(mem_0_144_W0_addr),
    .W0_clk(mem_0_144_W0_clk),
    .W0_data(mem_0_144_W0_data),
    .W0_en(mem_0_144_W0_en),
    .W0_mask(mem_0_144_W0_mask),
    .R0_addr(mem_0_144_R0_addr),
    .R0_clk(mem_0_144_R0_clk),
    .R0_data(mem_0_144_R0_data),
    .R0_en(mem_0_144_R0_en)
  );
  split_mem_0_ext mem_0_145 (
    .W0_addr(mem_0_145_W0_addr),
    .W0_clk(mem_0_145_W0_clk),
    .W0_data(mem_0_145_W0_data),
    .W0_en(mem_0_145_W0_en),
    .W0_mask(mem_0_145_W0_mask),
    .R0_addr(mem_0_145_R0_addr),
    .R0_clk(mem_0_145_R0_clk),
    .R0_data(mem_0_145_R0_data),
    .R0_en(mem_0_145_R0_en)
  );
  split_mem_0_ext mem_0_146 (
    .W0_addr(mem_0_146_W0_addr),
    .W0_clk(mem_0_146_W0_clk),
    .W0_data(mem_0_146_W0_data),
    .W0_en(mem_0_146_W0_en),
    .W0_mask(mem_0_146_W0_mask),
    .R0_addr(mem_0_146_R0_addr),
    .R0_clk(mem_0_146_R0_clk),
    .R0_data(mem_0_146_R0_data),
    .R0_en(mem_0_146_R0_en)
  );
  split_mem_0_ext mem_0_147 (
    .W0_addr(mem_0_147_W0_addr),
    .W0_clk(mem_0_147_W0_clk),
    .W0_data(mem_0_147_W0_data),
    .W0_en(mem_0_147_W0_en),
    .W0_mask(mem_0_147_W0_mask),
    .R0_addr(mem_0_147_R0_addr),
    .R0_clk(mem_0_147_R0_clk),
    .R0_data(mem_0_147_R0_data),
    .R0_en(mem_0_147_R0_en)
  );
  split_mem_0_ext mem_0_148 (
    .W0_addr(mem_0_148_W0_addr),
    .W0_clk(mem_0_148_W0_clk),
    .W0_data(mem_0_148_W0_data),
    .W0_en(mem_0_148_W0_en),
    .W0_mask(mem_0_148_W0_mask),
    .R0_addr(mem_0_148_R0_addr),
    .R0_clk(mem_0_148_R0_clk),
    .R0_data(mem_0_148_R0_data),
    .R0_en(mem_0_148_R0_en)
  );
  split_mem_0_ext mem_0_149 (
    .W0_addr(mem_0_149_W0_addr),
    .W0_clk(mem_0_149_W0_clk),
    .W0_data(mem_0_149_W0_data),
    .W0_en(mem_0_149_W0_en),
    .W0_mask(mem_0_149_W0_mask),
    .R0_addr(mem_0_149_R0_addr),
    .R0_clk(mem_0_149_R0_clk),
    .R0_data(mem_0_149_R0_data),
    .R0_en(mem_0_149_R0_en)
  );
  split_mem_0_ext mem_0_150 (
    .W0_addr(mem_0_150_W0_addr),
    .W0_clk(mem_0_150_W0_clk),
    .W0_data(mem_0_150_W0_data),
    .W0_en(mem_0_150_W0_en),
    .W0_mask(mem_0_150_W0_mask),
    .R0_addr(mem_0_150_R0_addr),
    .R0_clk(mem_0_150_R0_clk),
    .R0_data(mem_0_150_R0_data),
    .R0_en(mem_0_150_R0_en)
  );
  split_mem_0_ext mem_0_151 (
    .W0_addr(mem_0_151_W0_addr),
    .W0_clk(mem_0_151_W0_clk),
    .W0_data(mem_0_151_W0_data),
    .W0_en(mem_0_151_W0_en),
    .W0_mask(mem_0_151_W0_mask),
    .R0_addr(mem_0_151_R0_addr),
    .R0_clk(mem_0_151_R0_clk),
    .R0_data(mem_0_151_R0_data),
    .R0_en(mem_0_151_R0_en)
  );
  split_mem_0_ext mem_0_152 (
    .W0_addr(mem_0_152_W0_addr),
    .W0_clk(mem_0_152_W0_clk),
    .W0_data(mem_0_152_W0_data),
    .W0_en(mem_0_152_W0_en),
    .W0_mask(mem_0_152_W0_mask),
    .R0_addr(mem_0_152_R0_addr),
    .R0_clk(mem_0_152_R0_clk),
    .R0_data(mem_0_152_R0_data),
    .R0_en(mem_0_152_R0_en)
  );
  split_mem_0_ext mem_0_153 (
    .W0_addr(mem_0_153_W0_addr),
    .W0_clk(mem_0_153_W0_clk),
    .W0_data(mem_0_153_W0_data),
    .W0_en(mem_0_153_W0_en),
    .W0_mask(mem_0_153_W0_mask),
    .R0_addr(mem_0_153_R0_addr),
    .R0_clk(mem_0_153_R0_clk),
    .R0_data(mem_0_153_R0_data),
    .R0_en(mem_0_153_R0_en)
  );
  split_mem_0_ext mem_0_154 (
    .W0_addr(mem_0_154_W0_addr),
    .W0_clk(mem_0_154_W0_clk),
    .W0_data(mem_0_154_W0_data),
    .W0_en(mem_0_154_W0_en),
    .W0_mask(mem_0_154_W0_mask),
    .R0_addr(mem_0_154_R0_addr),
    .R0_clk(mem_0_154_R0_clk),
    .R0_data(mem_0_154_R0_data),
    .R0_en(mem_0_154_R0_en)
  );
  split_mem_0_ext mem_0_155 (
    .W0_addr(mem_0_155_W0_addr),
    .W0_clk(mem_0_155_W0_clk),
    .W0_data(mem_0_155_W0_data),
    .W0_en(mem_0_155_W0_en),
    .W0_mask(mem_0_155_W0_mask),
    .R0_addr(mem_0_155_R0_addr),
    .R0_clk(mem_0_155_R0_clk),
    .R0_data(mem_0_155_R0_data),
    .R0_en(mem_0_155_R0_en)
  );
  split_mem_0_ext mem_0_156 (
    .W0_addr(mem_0_156_W0_addr),
    .W0_clk(mem_0_156_W0_clk),
    .W0_data(mem_0_156_W0_data),
    .W0_en(mem_0_156_W0_en),
    .W0_mask(mem_0_156_W0_mask),
    .R0_addr(mem_0_156_R0_addr),
    .R0_clk(mem_0_156_R0_clk),
    .R0_data(mem_0_156_R0_data),
    .R0_en(mem_0_156_R0_en)
  );
  split_mem_0_ext mem_0_157 (
    .W0_addr(mem_0_157_W0_addr),
    .W0_clk(mem_0_157_W0_clk),
    .W0_data(mem_0_157_W0_data),
    .W0_en(mem_0_157_W0_en),
    .W0_mask(mem_0_157_W0_mask),
    .R0_addr(mem_0_157_R0_addr),
    .R0_clk(mem_0_157_R0_clk),
    .R0_data(mem_0_157_R0_data),
    .R0_en(mem_0_157_R0_en)
  );
  split_mem_0_ext mem_0_158 (
    .W0_addr(mem_0_158_W0_addr),
    .W0_clk(mem_0_158_W0_clk),
    .W0_data(mem_0_158_W0_data),
    .W0_en(mem_0_158_W0_en),
    .W0_mask(mem_0_158_W0_mask),
    .R0_addr(mem_0_158_R0_addr),
    .R0_clk(mem_0_158_R0_clk),
    .R0_data(mem_0_158_R0_data),
    .R0_en(mem_0_158_R0_en)
  );
  split_mem_0_ext mem_0_159 (
    .W0_addr(mem_0_159_W0_addr),
    .W0_clk(mem_0_159_W0_clk),
    .W0_data(mem_0_159_W0_data),
    .W0_en(mem_0_159_W0_en),
    .W0_mask(mem_0_159_W0_mask),
    .R0_addr(mem_0_159_R0_addr),
    .R0_clk(mem_0_159_R0_clk),
    .R0_data(mem_0_159_R0_data),
    .R0_en(mem_0_159_R0_en)
  );
  split_mem_0_ext mem_0_160 (
    .W0_addr(mem_0_160_W0_addr),
    .W0_clk(mem_0_160_W0_clk),
    .W0_data(mem_0_160_W0_data),
    .W0_en(mem_0_160_W0_en),
    .W0_mask(mem_0_160_W0_mask),
    .R0_addr(mem_0_160_R0_addr),
    .R0_clk(mem_0_160_R0_clk),
    .R0_data(mem_0_160_R0_data),
    .R0_en(mem_0_160_R0_en)
  );
  split_mem_0_ext mem_0_161 (
    .W0_addr(mem_0_161_W0_addr),
    .W0_clk(mem_0_161_W0_clk),
    .W0_data(mem_0_161_W0_data),
    .W0_en(mem_0_161_W0_en),
    .W0_mask(mem_0_161_W0_mask),
    .R0_addr(mem_0_161_R0_addr),
    .R0_clk(mem_0_161_R0_clk),
    .R0_data(mem_0_161_R0_data),
    .R0_en(mem_0_161_R0_en)
  );
  split_mem_0_ext mem_0_162 (
    .W0_addr(mem_0_162_W0_addr),
    .W0_clk(mem_0_162_W0_clk),
    .W0_data(mem_0_162_W0_data),
    .W0_en(mem_0_162_W0_en),
    .W0_mask(mem_0_162_W0_mask),
    .R0_addr(mem_0_162_R0_addr),
    .R0_clk(mem_0_162_R0_clk),
    .R0_data(mem_0_162_R0_data),
    .R0_en(mem_0_162_R0_en)
  );
  split_mem_0_ext mem_0_163 (
    .W0_addr(mem_0_163_W0_addr),
    .W0_clk(mem_0_163_W0_clk),
    .W0_data(mem_0_163_W0_data),
    .W0_en(mem_0_163_W0_en),
    .W0_mask(mem_0_163_W0_mask),
    .R0_addr(mem_0_163_R0_addr),
    .R0_clk(mem_0_163_R0_clk),
    .R0_data(mem_0_163_R0_data),
    .R0_en(mem_0_163_R0_en)
  );
  split_mem_0_ext mem_0_164 (
    .W0_addr(mem_0_164_W0_addr),
    .W0_clk(mem_0_164_W0_clk),
    .W0_data(mem_0_164_W0_data),
    .W0_en(mem_0_164_W0_en),
    .W0_mask(mem_0_164_W0_mask),
    .R0_addr(mem_0_164_R0_addr),
    .R0_clk(mem_0_164_R0_clk),
    .R0_data(mem_0_164_R0_data),
    .R0_en(mem_0_164_R0_en)
  );
  split_mem_0_ext mem_0_165 (
    .W0_addr(mem_0_165_W0_addr),
    .W0_clk(mem_0_165_W0_clk),
    .W0_data(mem_0_165_W0_data),
    .W0_en(mem_0_165_W0_en),
    .W0_mask(mem_0_165_W0_mask),
    .R0_addr(mem_0_165_R0_addr),
    .R0_clk(mem_0_165_R0_clk),
    .R0_data(mem_0_165_R0_data),
    .R0_en(mem_0_165_R0_en)
  );
  split_mem_0_ext mem_0_166 (
    .W0_addr(mem_0_166_W0_addr),
    .W0_clk(mem_0_166_W0_clk),
    .W0_data(mem_0_166_W0_data),
    .W0_en(mem_0_166_W0_en),
    .W0_mask(mem_0_166_W0_mask),
    .R0_addr(mem_0_166_R0_addr),
    .R0_clk(mem_0_166_R0_clk),
    .R0_data(mem_0_166_R0_data),
    .R0_en(mem_0_166_R0_en)
  );
  split_mem_0_ext mem_0_167 (
    .W0_addr(mem_0_167_W0_addr),
    .W0_clk(mem_0_167_W0_clk),
    .W0_data(mem_0_167_W0_data),
    .W0_en(mem_0_167_W0_en),
    .W0_mask(mem_0_167_W0_mask),
    .R0_addr(mem_0_167_R0_addr),
    .R0_clk(mem_0_167_R0_clk),
    .R0_data(mem_0_167_R0_data),
    .R0_en(mem_0_167_R0_en)
  );
  split_mem_0_ext mem_0_168 (
    .W0_addr(mem_0_168_W0_addr),
    .W0_clk(mem_0_168_W0_clk),
    .W0_data(mem_0_168_W0_data),
    .W0_en(mem_0_168_W0_en),
    .W0_mask(mem_0_168_W0_mask),
    .R0_addr(mem_0_168_R0_addr),
    .R0_clk(mem_0_168_R0_clk),
    .R0_data(mem_0_168_R0_data),
    .R0_en(mem_0_168_R0_en)
  );
  split_mem_0_ext mem_0_169 (
    .W0_addr(mem_0_169_W0_addr),
    .W0_clk(mem_0_169_W0_clk),
    .W0_data(mem_0_169_W0_data),
    .W0_en(mem_0_169_W0_en),
    .W0_mask(mem_0_169_W0_mask),
    .R0_addr(mem_0_169_R0_addr),
    .R0_clk(mem_0_169_R0_clk),
    .R0_data(mem_0_169_R0_data),
    .R0_en(mem_0_169_R0_en)
  );
  split_mem_0_ext mem_0_170 (
    .W0_addr(mem_0_170_W0_addr),
    .W0_clk(mem_0_170_W0_clk),
    .W0_data(mem_0_170_W0_data),
    .W0_en(mem_0_170_W0_en),
    .W0_mask(mem_0_170_W0_mask),
    .R0_addr(mem_0_170_R0_addr),
    .R0_clk(mem_0_170_R0_clk),
    .R0_data(mem_0_170_R0_data),
    .R0_en(mem_0_170_R0_en)
  );
  split_mem_0_ext mem_0_171 (
    .W0_addr(mem_0_171_W0_addr),
    .W0_clk(mem_0_171_W0_clk),
    .W0_data(mem_0_171_W0_data),
    .W0_en(mem_0_171_W0_en),
    .W0_mask(mem_0_171_W0_mask),
    .R0_addr(mem_0_171_R0_addr),
    .R0_clk(mem_0_171_R0_clk),
    .R0_data(mem_0_171_R0_data),
    .R0_en(mem_0_171_R0_en)
  );
  split_mem_0_ext mem_0_172 (
    .W0_addr(mem_0_172_W0_addr),
    .W0_clk(mem_0_172_W0_clk),
    .W0_data(mem_0_172_W0_data),
    .W0_en(mem_0_172_W0_en),
    .W0_mask(mem_0_172_W0_mask),
    .R0_addr(mem_0_172_R0_addr),
    .R0_clk(mem_0_172_R0_clk),
    .R0_data(mem_0_172_R0_data),
    .R0_en(mem_0_172_R0_en)
  );
  split_mem_0_ext mem_0_173 (
    .W0_addr(mem_0_173_W0_addr),
    .W0_clk(mem_0_173_W0_clk),
    .W0_data(mem_0_173_W0_data),
    .W0_en(mem_0_173_W0_en),
    .W0_mask(mem_0_173_W0_mask),
    .R0_addr(mem_0_173_R0_addr),
    .R0_clk(mem_0_173_R0_clk),
    .R0_data(mem_0_173_R0_data),
    .R0_en(mem_0_173_R0_en)
  );
  split_mem_0_ext mem_0_174 (
    .W0_addr(mem_0_174_W0_addr),
    .W0_clk(mem_0_174_W0_clk),
    .W0_data(mem_0_174_W0_data),
    .W0_en(mem_0_174_W0_en),
    .W0_mask(mem_0_174_W0_mask),
    .R0_addr(mem_0_174_R0_addr),
    .R0_clk(mem_0_174_R0_clk),
    .R0_data(mem_0_174_R0_data),
    .R0_en(mem_0_174_R0_en)
  );
  split_mem_0_ext mem_0_175 (
    .W0_addr(mem_0_175_W0_addr),
    .W0_clk(mem_0_175_W0_clk),
    .W0_data(mem_0_175_W0_data),
    .W0_en(mem_0_175_W0_en),
    .W0_mask(mem_0_175_W0_mask),
    .R0_addr(mem_0_175_R0_addr),
    .R0_clk(mem_0_175_R0_clk),
    .R0_data(mem_0_175_R0_data),
    .R0_en(mem_0_175_R0_en)
  );
  split_mem_0_ext mem_0_176 (
    .W0_addr(mem_0_176_W0_addr),
    .W0_clk(mem_0_176_W0_clk),
    .W0_data(mem_0_176_W0_data),
    .W0_en(mem_0_176_W0_en),
    .W0_mask(mem_0_176_W0_mask),
    .R0_addr(mem_0_176_R0_addr),
    .R0_clk(mem_0_176_R0_clk),
    .R0_data(mem_0_176_R0_data),
    .R0_en(mem_0_176_R0_en)
  );
  split_mem_0_ext mem_0_177 (
    .W0_addr(mem_0_177_W0_addr),
    .W0_clk(mem_0_177_W0_clk),
    .W0_data(mem_0_177_W0_data),
    .W0_en(mem_0_177_W0_en),
    .W0_mask(mem_0_177_W0_mask),
    .R0_addr(mem_0_177_R0_addr),
    .R0_clk(mem_0_177_R0_clk),
    .R0_data(mem_0_177_R0_data),
    .R0_en(mem_0_177_R0_en)
  );
  split_mem_0_ext mem_0_178 (
    .W0_addr(mem_0_178_W0_addr),
    .W0_clk(mem_0_178_W0_clk),
    .W0_data(mem_0_178_W0_data),
    .W0_en(mem_0_178_W0_en),
    .W0_mask(mem_0_178_W0_mask),
    .R0_addr(mem_0_178_R0_addr),
    .R0_clk(mem_0_178_R0_clk),
    .R0_data(mem_0_178_R0_data),
    .R0_en(mem_0_178_R0_en)
  );
  split_mem_0_ext mem_0_179 (
    .W0_addr(mem_0_179_W0_addr),
    .W0_clk(mem_0_179_W0_clk),
    .W0_data(mem_0_179_W0_data),
    .W0_en(mem_0_179_W0_en),
    .W0_mask(mem_0_179_W0_mask),
    .R0_addr(mem_0_179_R0_addr),
    .R0_clk(mem_0_179_R0_clk),
    .R0_data(mem_0_179_R0_data),
    .R0_en(mem_0_179_R0_en)
  );
  split_mem_0_ext mem_0_180 (
    .W0_addr(mem_0_180_W0_addr),
    .W0_clk(mem_0_180_W0_clk),
    .W0_data(mem_0_180_W0_data),
    .W0_en(mem_0_180_W0_en),
    .W0_mask(mem_0_180_W0_mask),
    .R0_addr(mem_0_180_R0_addr),
    .R0_clk(mem_0_180_R0_clk),
    .R0_data(mem_0_180_R0_data),
    .R0_en(mem_0_180_R0_en)
  );
  split_mem_0_ext mem_0_181 (
    .W0_addr(mem_0_181_W0_addr),
    .W0_clk(mem_0_181_W0_clk),
    .W0_data(mem_0_181_W0_data),
    .W0_en(mem_0_181_W0_en),
    .W0_mask(mem_0_181_W0_mask),
    .R0_addr(mem_0_181_R0_addr),
    .R0_clk(mem_0_181_R0_clk),
    .R0_data(mem_0_181_R0_data),
    .R0_en(mem_0_181_R0_en)
  );
  split_mem_0_ext mem_0_182 (
    .W0_addr(mem_0_182_W0_addr),
    .W0_clk(mem_0_182_W0_clk),
    .W0_data(mem_0_182_W0_data),
    .W0_en(mem_0_182_W0_en),
    .W0_mask(mem_0_182_W0_mask),
    .R0_addr(mem_0_182_R0_addr),
    .R0_clk(mem_0_182_R0_clk),
    .R0_data(mem_0_182_R0_data),
    .R0_en(mem_0_182_R0_en)
  );
  split_mem_0_ext mem_0_183 (
    .W0_addr(mem_0_183_W0_addr),
    .W0_clk(mem_0_183_W0_clk),
    .W0_data(mem_0_183_W0_data),
    .W0_en(mem_0_183_W0_en),
    .W0_mask(mem_0_183_W0_mask),
    .R0_addr(mem_0_183_R0_addr),
    .R0_clk(mem_0_183_R0_clk),
    .R0_data(mem_0_183_R0_data),
    .R0_en(mem_0_183_R0_en)
  );
  split_mem_0_ext mem_0_184 (
    .W0_addr(mem_0_184_W0_addr),
    .W0_clk(mem_0_184_W0_clk),
    .W0_data(mem_0_184_W0_data),
    .W0_en(mem_0_184_W0_en),
    .W0_mask(mem_0_184_W0_mask),
    .R0_addr(mem_0_184_R0_addr),
    .R0_clk(mem_0_184_R0_clk),
    .R0_data(mem_0_184_R0_data),
    .R0_en(mem_0_184_R0_en)
  );
  split_mem_0_ext mem_0_185 (
    .W0_addr(mem_0_185_W0_addr),
    .W0_clk(mem_0_185_W0_clk),
    .W0_data(mem_0_185_W0_data),
    .W0_en(mem_0_185_W0_en),
    .W0_mask(mem_0_185_W0_mask),
    .R0_addr(mem_0_185_R0_addr),
    .R0_clk(mem_0_185_R0_clk),
    .R0_data(mem_0_185_R0_data),
    .R0_en(mem_0_185_R0_en)
  );
  split_mem_0_ext mem_0_186 (
    .W0_addr(mem_0_186_W0_addr),
    .W0_clk(mem_0_186_W0_clk),
    .W0_data(mem_0_186_W0_data),
    .W0_en(mem_0_186_W0_en),
    .W0_mask(mem_0_186_W0_mask),
    .R0_addr(mem_0_186_R0_addr),
    .R0_clk(mem_0_186_R0_clk),
    .R0_data(mem_0_186_R0_data),
    .R0_en(mem_0_186_R0_en)
  );
  split_mem_0_ext mem_0_187 (
    .W0_addr(mem_0_187_W0_addr),
    .W0_clk(mem_0_187_W0_clk),
    .W0_data(mem_0_187_W0_data),
    .W0_en(mem_0_187_W0_en),
    .W0_mask(mem_0_187_W0_mask),
    .R0_addr(mem_0_187_R0_addr),
    .R0_clk(mem_0_187_R0_clk),
    .R0_data(mem_0_187_R0_data),
    .R0_en(mem_0_187_R0_en)
  );
  split_mem_0_ext mem_0_188 (
    .W0_addr(mem_0_188_W0_addr),
    .W0_clk(mem_0_188_W0_clk),
    .W0_data(mem_0_188_W0_data),
    .W0_en(mem_0_188_W0_en),
    .W0_mask(mem_0_188_W0_mask),
    .R0_addr(mem_0_188_R0_addr),
    .R0_clk(mem_0_188_R0_clk),
    .R0_data(mem_0_188_R0_data),
    .R0_en(mem_0_188_R0_en)
  );
  split_mem_0_ext mem_0_189 (
    .W0_addr(mem_0_189_W0_addr),
    .W0_clk(mem_0_189_W0_clk),
    .W0_data(mem_0_189_W0_data),
    .W0_en(mem_0_189_W0_en),
    .W0_mask(mem_0_189_W0_mask),
    .R0_addr(mem_0_189_R0_addr),
    .R0_clk(mem_0_189_R0_clk),
    .R0_data(mem_0_189_R0_data),
    .R0_en(mem_0_189_R0_en)
  );
  split_mem_0_ext mem_0_190 (
    .W0_addr(mem_0_190_W0_addr),
    .W0_clk(mem_0_190_W0_clk),
    .W0_data(mem_0_190_W0_data),
    .W0_en(mem_0_190_W0_en),
    .W0_mask(mem_0_190_W0_mask),
    .R0_addr(mem_0_190_R0_addr),
    .R0_clk(mem_0_190_R0_clk),
    .R0_data(mem_0_190_R0_data),
    .R0_en(mem_0_190_R0_en)
  );
  split_mem_0_ext mem_0_191 (
    .W0_addr(mem_0_191_W0_addr),
    .W0_clk(mem_0_191_W0_clk),
    .W0_data(mem_0_191_W0_data),
    .W0_en(mem_0_191_W0_en),
    .W0_mask(mem_0_191_W0_mask),
    .R0_addr(mem_0_191_R0_addr),
    .R0_clk(mem_0_191_R0_clk),
    .R0_data(mem_0_191_R0_data),
    .R0_en(mem_0_191_R0_en)
  );
  split_mem_0_ext mem_0_192 (
    .W0_addr(mem_0_192_W0_addr),
    .W0_clk(mem_0_192_W0_clk),
    .W0_data(mem_0_192_W0_data),
    .W0_en(mem_0_192_W0_en),
    .W0_mask(mem_0_192_W0_mask),
    .R0_addr(mem_0_192_R0_addr),
    .R0_clk(mem_0_192_R0_clk),
    .R0_data(mem_0_192_R0_data),
    .R0_en(mem_0_192_R0_en)
  );
  split_mem_0_ext mem_0_193 (
    .W0_addr(mem_0_193_W0_addr),
    .W0_clk(mem_0_193_W0_clk),
    .W0_data(mem_0_193_W0_data),
    .W0_en(mem_0_193_W0_en),
    .W0_mask(mem_0_193_W0_mask),
    .R0_addr(mem_0_193_R0_addr),
    .R0_clk(mem_0_193_R0_clk),
    .R0_data(mem_0_193_R0_data),
    .R0_en(mem_0_193_R0_en)
  );
  split_mem_0_ext mem_0_194 (
    .W0_addr(mem_0_194_W0_addr),
    .W0_clk(mem_0_194_W0_clk),
    .W0_data(mem_0_194_W0_data),
    .W0_en(mem_0_194_W0_en),
    .W0_mask(mem_0_194_W0_mask),
    .R0_addr(mem_0_194_R0_addr),
    .R0_clk(mem_0_194_R0_clk),
    .R0_data(mem_0_194_R0_data),
    .R0_en(mem_0_194_R0_en)
  );
  split_mem_0_ext mem_0_195 (
    .W0_addr(mem_0_195_W0_addr),
    .W0_clk(mem_0_195_W0_clk),
    .W0_data(mem_0_195_W0_data),
    .W0_en(mem_0_195_W0_en),
    .W0_mask(mem_0_195_W0_mask),
    .R0_addr(mem_0_195_R0_addr),
    .R0_clk(mem_0_195_R0_clk),
    .R0_data(mem_0_195_R0_data),
    .R0_en(mem_0_195_R0_en)
  );
  split_mem_0_ext mem_0_196 (
    .W0_addr(mem_0_196_W0_addr),
    .W0_clk(mem_0_196_W0_clk),
    .W0_data(mem_0_196_W0_data),
    .W0_en(mem_0_196_W0_en),
    .W0_mask(mem_0_196_W0_mask),
    .R0_addr(mem_0_196_R0_addr),
    .R0_clk(mem_0_196_R0_clk),
    .R0_data(mem_0_196_R0_data),
    .R0_en(mem_0_196_R0_en)
  );
  split_mem_0_ext mem_0_197 (
    .W0_addr(mem_0_197_W0_addr),
    .W0_clk(mem_0_197_W0_clk),
    .W0_data(mem_0_197_W0_data),
    .W0_en(mem_0_197_W0_en),
    .W0_mask(mem_0_197_W0_mask),
    .R0_addr(mem_0_197_R0_addr),
    .R0_clk(mem_0_197_R0_clk),
    .R0_data(mem_0_197_R0_data),
    .R0_en(mem_0_197_R0_en)
  );
  split_mem_0_ext mem_0_198 (
    .W0_addr(mem_0_198_W0_addr),
    .W0_clk(mem_0_198_W0_clk),
    .W0_data(mem_0_198_W0_data),
    .W0_en(mem_0_198_W0_en),
    .W0_mask(mem_0_198_W0_mask),
    .R0_addr(mem_0_198_R0_addr),
    .R0_clk(mem_0_198_R0_clk),
    .R0_data(mem_0_198_R0_data),
    .R0_en(mem_0_198_R0_en)
  );
  split_mem_0_ext mem_0_199 (
    .W0_addr(mem_0_199_W0_addr),
    .W0_clk(mem_0_199_W0_clk),
    .W0_data(mem_0_199_W0_data),
    .W0_en(mem_0_199_W0_en),
    .W0_mask(mem_0_199_W0_mask),
    .R0_addr(mem_0_199_R0_addr),
    .R0_clk(mem_0_199_R0_clk),
    .R0_data(mem_0_199_R0_data),
    .R0_en(mem_0_199_R0_en)
  );
  split_mem_0_ext mem_0_200 (
    .W0_addr(mem_0_200_W0_addr),
    .W0_clk(mem_0_200_W0_clk),
    .W0_data(mem_0_200_W0_data),
    .W0_en(mem_0_200_W0_en),
    .W0_mask(mem_0_200_W0_mask),
    .R0_addr(mem_0_200_R0_addr),
    .R0_clk(mem_0_200_R0_clk),
    .R0_data(mem_0_200_R0_data),
    .R0_en(mem_0_200_R0_en)
  );
  split_mem_0_ext mem_0_201 (
    .W0_addr(mem_0_201_W0_addr),
    .W0_clk(mem_0_201_W0_clk),
    .W0_data(mem_0_201_W0_data),
    .W0_en(mem_0_201_W0_en),
    .W0_mask(mem_0_201_W0_mask),
    .R0_addr(mem_0_201_R0_addr),
    .R0_clk(mem_0_201_R0_clk),
    .R0_data(mem_0_201_R0_data),
    .R0_en(mem_0_201_R0_en)
  );
  split_mem_0_ext mem_0_202 (
    .W0_addr(mem_0_202_W0_addr),
    .W0_clk(mem_0_202_W0_clk),
    .W0_data(mem_0_202_W0_data),
    .W0_en(mem_0_202_W0_en),
    .W0_mask(mem_0_202_W0_mask),
    .R0_addr(mem_0_202_R0_addr),
    .R0_clk(mem_0_202_R0_clk),
    .R0_data(mem_0_202_R0_data),
    .R0_en(mem_0_202_R0_en)
  );
  split_mem_0_ext mem_0_203 (
    .W0_addr(mem_0_203_W0_addr),
    .W0_clk(mem_0_203_W0_clk),
    .W0_data(mem_0_203_W0_data),
    .W0_en(mem_0_203_W0_en),
    .W0_mask(mem_0_203_W0_mask),
    .R0_addr(mem_0_203_R0_addr),
    .R0_clk(mem_0_203_R0_clk),
    .R0_data(mem_0_203_R0_data),
    .R0_en(mem_0_203_R0_en)
  );
  split_mem_0_ext mem_0_204 (
    .W0_addr(mem_0_204_W0_addr),
    .W0_clk(mem_0_204_W0_clk),
    .W0_data(mem_0_204_W0_data),
    .W0_en(mem_0_204_W0_en),
    .W0_mask(mem_0_204_W0_mask),
    .R0_addr(mem_0_204_R0_addr),
    .R0_clk(mem_0_204_R0_clk),
    .R0_data(mem_0_204_R0_data),
    .R0_en(mem_0_204_R0_en)
  );
  split_mem_0_ext mem_0_205 (
    .W0_addr(mem_0_205_W0_addr),
    .W0_clk(mem_0_205_W0_clk),
    .W0_data(mem_0_205_W0_data),
    .W0_en(mem_0_205_W0_en),
    .W0_mask(mem_0_205_W0_mask),
    .R0_addr(mem_0_205_R0_addr),
    .R0_clk(mem_0_205_R0_clk),
    .R0_data(mem_0_205_R0_data),
    .R0_en(mem_0_205_R0_en)
  );
  split_mem_0_ext mem_0_206 (
    .W0_addr(mem_0_206_W0_addr),
    .W0_clk(mem_0_206_W0_clk),
    .W0_data(mem_0_206_W0_data),
    .W0_en(mem_0_206_W0_en),
    .W0_mask(mem_0_206_W0_mask),
    .R0_addr(mem_0_206_R0_addr),
    .R0_clk(mem_0_206_R0_clk),
    .R0_data(mem_0_206_R0_data),
    .R0_en(mem_0_206_R0_en)
  );
  split_mem_0_ext mem_0_207 (
    .W0_addr(mem_0_207_W0_addr),
    .W0_clk(mem_0_207_W0_clk),
    .W0_data(mem_0_207_W0_data),
    .W0_en(mem_0_207_W0_en),
    .W0_mask(mem_0_207_W0_mask),
    .R0_addr(mem_0_207_R0_addr),
    .R0_clk(mem_0_207_R0_clk),
    .R0_data(mem_0_207_R0_data),
    .R0_en(mem_0_207_R0_en)
  );
  split_mem_0_ext mem_0_208 (
    .W0_addr(mem_0_208_W0_addr),
    .W0_clk(mem_0_208_W0_clk),
    .W0_data(mem_0_208_W0_data),
    .W0_en(mem_0_208_W0_en),
    .W0_mask(mem_0_208_W0_mask),
    .R0_addr(mem_0_208_R0_addr),
    .R0_clk(mem_0_208_R0_clk),
    .R0_data(mem_0_208_R0_data),
    .R0_en(mem_0_208_R0_en)
  );
  split_mem_0_ext mem_0_209 (
    .W0_addr(mem_0_209_W0_addr),
    .W0_clk(mem_0_209_W0_clk),
    .W0_data(mem_0_209_W0_data),
    .W0_en(mem_0_209_W0_en),
    .W0_mask(mem_0_209_W0_mask),
    .R0_addr(mem_0_209_R0_addr),
    .R0_clk(mem_0_209_R0_clk),
    .R0_data(mem_0_209_R0_data),
    .R0_en(mem_0_209_R0_en)
  );
  split_mem_0_ext mem_0_210 (
    .W0_addr(mem_0_210_W0_addr),
    .W0_clk(mem_0_210_W0_clk),
    .W0_data(mem_0_210_W0_data),
    .W0_en(mem_0_210_W0_en),
    .W0_mask(mem_0_210_W0_mask),
    .R0_addr(mem_0_210_R0_addr),
    .R0_clk(mem_0_210_R0_clk),
    .R0_data(mem_0_210_R0_data),
    .R0_en(mem_0_210_R0_en)
  );
  split_mem_0_ext mem_0_211 (
    .W0_addr(mem_0_211_W0_addr),
    .W0_clk(mem_0_211_W0_clk),
    .W0_data(mem_0_211_W0_data),
    .W0_en(mem_0_211_W0_en),
    .W0_mask(mem_0_211_W0_mask),
    .R0_addr(mem_0_211_R0_addr),
    .R0_clk(mem_0_211_R0_clk),
    .R0_data(mem_0_211_R0_data),
    .R0_en(mem_0_211_R0_en)
  );
  split_mem_0_ext mem_0_212 (
    .W0_addr(mem_0_212_W0_addr),
    .W0_clk(mem_0_212_W0_clk),
    .W0_data(mem_0_212_W0_data),
    .W0_en(mem_0_212_W0_en),
    .W0_mask(mem_0_212_W0_mask),
    .R0_addr(mem_0_212_R0_addr),
    .R0_clk(mem_0_212_R0_clk),
    .R0_data(mem_0_212_R0_data),
    .R0_en(mem_0_212_R0_en)
  );
  split_mem_0_ext mem_0_213 (
    .W0_addr(mem_0_213_W0_addr),
    .W0_clk(mem_0_213_W0_clk),
    .W0_data(mem_0_213_W0_data),
    .W0_en(mem_0_213_W0_en),
    .W0_mask(mem_0_213_W0_mask),
    .R0_addr(mem_0_213_R0_addr),
    .R0_clk(mem_0_213_R0_clk),
    .R0_data(mem_0_213_R0_data),
    .R0_en(mem_0_213_R0_en)
  );
  split_mem_0_ext mem_0_214 (
    .W0_addr(mem_0_214_W0_addr),
    .W0_clk(mem_0_214_W0_clk),
    .W0_data(mem_0_214_W0_data),
    .W0_en(mem_0_214_W0_en),
    .W0_mask(mem_0_214_W0_mask),
    .R0_addr(mem_0_214_R0_addr),
    .R0_clk(mem_0_214_R0_clk),
    .R0_data(mem_0_214_R0_data),
    .R0_en(mem_0_214_R0_en)
  );
  split_mem_0_ext mem_0_215 (
    .W0_addr(mem_0_215_W0_addr),
    .W0_clk(mem_0_215_W0_clk),
    .W0_data(mem_0_215_W0_data),
    .W0_en(mem_0_215_W0_en),
    .W0_mask(mem_0_215_W0_mask),
    .R0_addr(mem_0_215_R0_addr),
    .R0_clk(mem_0_215_R0_clk),
    .R0_data(mem_0_215_R0_data),
    .R0_en(mem_0_215_R0_en)
  );
  split_mem_0_ext mem_0_216 (
    .W0_addr(mem_0_216_W0_addr),
    .W0_clk(mem_0_216_W0_clk),
    .W0_data(mem_0_216_W0_data),
    .W0_en(mem_0_216_W0_en),
    .W0_mask(mem_0_216_W0_mask),
    .R0_addr(mem_0_216_R0_addr),
    .R0_clk(mem_0_216_R0_clk),
    .R0_data(mem_0_216_R0_data),
    .R0_en(mem_0_216_R0_en)
  );
  split_mem_0_ext mem_0_217 (
    .W0_addr(mem_0_217_W0_addr),
    .W0_clk(mem_0_217_W0_clk),
    .W0_data(mem_0_217_W0_data),
    .W0_en(mem_0_217_W0_en),
    .W0_mask(mem_0_217_W0_mask),
    .R0_addr(mem_0_217_R0_addr),
    .R0_clk(mem_0_217_R0_clk),
    .R0_data(mem_0_217_R0_data),
    .R0_en(mem_0_217_R0_en)
  );
  split_mem_0_ext mem_0_218 (
    .W0_addr(mem_0_218_W0_addr),
    .W0_clk(mem_0_218_W0_clk),
    .W0_data(mem_0_218_W0_data),
    .W0_en(mem_0_218_W0_en),
    .W0_mask(mem_0_218_W0_mask),
    .R0_addr(mem_0_218_R0_addr),
    .R0_clk(mem_0_218_R0_clk),
    .R0_data(mem_0_218_R0_data),
    .R0_en(mem_0_218_R0_en)
  );
  split_mem_0_ext mem_0_219 (
    .W0_addr(mem_0_219_W0_addr),
    .W0_clk(mem_0_219_W0_clk),
    .W0_data(mem_0_219_W0_data),
    .W0_en(mem_0_219_W0_en),
    .W0_mask(mem_0_219_W0_mask),
    .R0_addr(mem_0_219_R0_addr),
    .R0_clk(mem_0_219_R0_clk),
    .R0_data(mem_0_219_R0_data),
    .R0_en(mem_0_219_R0_en)
  );
  split_mem_0_ext mem_0_220 (
    .W0_addr(mem_0_220_W0_addr),
    .W0_clk(mem_0_220_W0_clk),
    .W0_data(mem_0_220_W0_data),
    .W0_en(mem_0_220_W0_en),
    .W0_mask(mem_0_220_W0_mask),
    .R0_addr(mem_0_220_R0_addr),
    .R0_clk(mem_0_220_R0_clk),
    .R0_data(mem_0_220_R0_data),
    .R0_en(mem_0_220_R0_en)
  );
  split_mem_0_ext mem_0_221 (
    .W0_addr(mem_0_221_W0_addr),
    .W0_clk(mem_0_221_W0_clk),
    .W0_data(mem_0_221_W0_data),
    .W0_en(mem_0_221_W0_en),
    .W0_mask(mem_0_221_W0_mask),
    .R0_addr(mem_0_221_R0_addr),
    .R0_clk(mem_0_221_R0_clk),
    .R0_data(mem_0_221_R0_data),
    .R0_en(mem_0_221_R0_en)
  );
  split_mem_0_ext mem_0_222 (
    .W0_addr(mem_0_222_W0_addr),
    .W0_clk(mem_0_222_W0_clk),
    .W0_data(mem_0_222_W0_data),
    .W0_en(mem_0_222_W0_en),
    .W0_mask(mem_0_222_W0_mask),
    .R0_addr(mem_0_222_R0_addr),
    .R0_clk(mem_0_222_R0_clk),
    .R0_data(mem_0_222_R0_data),
    .R0_en(mem_0_222_R0_en)
  );
  split_mem_0_ext mem_0_223 (
    .W0_addr(mem_0_223_W0_addr),
    .W0_clk(mem_0_223_W0_clk),
    .W0_data(mem_0_223_W0_data),
    .W0_en(mem_0_223_W0_en),
    .W0_mask(mem_0_223_W0_mask),
    .R0_addr(mem_0_223_R0_addr),
    .R0_clk(mem_0_223_R0_clk),
    .R0_data(mem_0_223_R0_data),
    .R0_en(mem_0_223_R0_en)
  );
  split_mem_0_ext mem_0_224 (
    .W0_addr(mem_0_224_W0_addr),
    .W0_clk(mem_0_224_W0_clk),
    .W0_data(mem_0_224_W0_data),
    .W0_en(mem_0_224_W0_en),
    .W0_mask(mem_0_224_W0_mask),
    .R0_addr(mem_0_224_R0_addr),
    .R0_clk(mem_0_224_R0_clk),
    .R0_data(mem_0_224_R0_data),
    .R0_en(mem_0_224_R0_en)
  );
  split_mem_0_ext mem_0_225 (
    .W0_addr(mem_0_225_W0_addr),
    .W0_clk(mem_0_225_W0_clk),
    .W0_data(mem_0_225_W0_data),
    .W0_en(mem_0_225_W0_en),
    .W0_mask(mem_0_225_W0_mask),
    .R0_addr(mem_0_225_R0_addr),
    .R0_clk(mem_0_225_R0_clk),
    .R0_data(mem_0_225_R0_data),
    .R0_en(mem_0_225_R0_en)
  );
  split_mem_0_ext mem_0_226 (
    .W0_addr(mem_0_226_W0_addr),
    .W0_clk(mem_0_226_W0_clk),
    .W0_data(mem_0_226_W0_data),
    .W0_en(mem_0_226_W0_en),
    .W0_mask(mem_0_226_W0_mask),
    .R0_addr(mem_0_226_R0_addr),
    .R0_clk(mem_0_226_R0_clk),
    .R0_data(mem_0_226_R0_data),
    .R0_en(mem_0_226_R0_en)
  );
  split_mem_0_ext mem_0_227 (
    .W0_addr(mem_0_227_W0_addr),
    .W0_clk(mem_0_227_W0_clk),
    .W0_data(mem_0_227_W0_data),
    .W0_en(mem_0_227_W0_en),
    .W0_mask(mem_0_227_W0_mask),
    .R0_addr(mem_0_227_R0_addr),
    .R0_clk(mem_0_227_R0_clk),
    .R0_data(mem_0_227_R0_data),
    .R0_en(mem_0_227_R0_en)
  );
  split_mem_0_ext mem_0_228 (
    .W0_addr(mem_0_228_W0_addr),
    .W0_clk(mem_0_228_W0_clk),
    .W0_data(mem_0_228_W0_data),
    .W0_en(mem_0_228_W0_en),
    .W0_mask(mem_0_228_W0_mask),
    .R0_addr(mem_0_228_R0_addr),
    .R0_clk(mem_0_228_R0_clk),
    .R0_data(mem_0_228_R0_data),
    .R0_en(mem_0_228_R0_en)
  );
  split_mem_0_ext mem_0_229 (
    .W0_addr(mem_0_229_W0_addr),
    .W0_clk(mem_0_229_W0_clk),
    .W0_data(mem_0_229_W0_data),
    .W0_en(mem_0_229_W0_en),
    .W0_mask(mem_0_229_W0_mask),
    .R0_addr(mem_0_229_R0_addr),
    .R0_clk(mem_0_229_R0_clk),
    .R0_data(mem_0_229_R0_data),
    .R0_en(mem_0_229_R0_en)
  );
  split_mem_0_ext mem_0_230 (
    .W0_addr(mem_0_230_W0_addr),
    .W0_clk(mem_0_230_W0_clk),
    .W0_data(mem_0_230_W0_data),
    .W0_en(mem_0_230_W0_en),
    .W0_mask(mem_0_230_W0_mask),
    .R0_addr(mem_0_230_R0_addr),
    .R0_clk(mem_0_230_R0_clk),
    .R0_data(mem_0_230_R0_data),
    .R0_en(mem_0_230_R0_en)
  );
  split_mem_0_ext mem_0_231 (
    .W0_addr(mem_0_231_W0_addr),
    .W0_clk(mem_0_231_W0_clk),
    .W0_data(mem_0_231_W0_data),
    .W0_en(mem_0_231_W0_en),
    .W0_mask(mem_0_231_W0_mask),
    .R0_addr(mem_0_231_R0_addr),
    .R0_clk(mem_0_231_R0_clk),
    .R0_data(mem_0_231_R0_data),
    .R0_en(mem_0_231_R0_en)
  );
  split_mem_0_ext mem_0_232 (
    .W0_addr(mem_0_232_W0_addr),
    .W0_clk(mem_0_232_W0_clk),
    .W0_data(mem_0_232_W0_data),
    .W0_en(mem_0_232_W0_en),
    .W0_mask(mem_0_232_W0_mask),
    .R0_addr(mem_0_232_R0_addr),
    .R0_clk(mem_0_232_R0_clk),
    .R0_data(mem_0_232_R0_data),
    .R0_en(mem_0_232_R0_en)
  );
  split_mem_0_ext mem_0_233 (
    .W0_addr(mem_0_233_W0_addr),
    .W0_clk(mem_0_233_W0_clk),
    .W0_data(mem_0_233_W0_data),
    .W0_en(mem_0_233_W0_en),
    .W0_mask(mem_0_233_W0_mask),
    .R0_addr(mem_0_233_R0_addr),
    .R0_clk(mem_0_233_R0_clk),
    .R0_data(mem_0_233_R0_data),
    .R0_en(mem_0_233_R0_en)
  );
  split_mem_0_ext mem_0_234 (
    .W0_addr(mem_0_234_W0_addr),
    .W0_clk(mem_0_234_W0_clk),
    .W0_data(mem_0_234_W0_data),
    .W0_en(mem_0_234_W0_en),
    .W0_mask(mem_0_234_W0_mask),
    .R0_addr(mem_0_234_R0_addr),
    .R0_clk(mem_0_234_R0_clk),
    .R0_data(mem_0_234_R0_data),
    .R0_en(mem_0_234_R0_en)
  );
  split_mem_0_ext mem_0_235 (
    .W0_addr(mem_0_235_W0_addr),
    .W0_clk(mem_0_235_W0_clk),
    .W0_data(mem_0_235_W0_data),
    .W0_en(mem_0_235_W0_en),
    .W0_mask(mem_0_235_W0_mask),
    .R0_addr(mem_0_235_R0_addr),
    .R0_clk(mem_0_235_R0_clk),
    .R0_data(mem_0_235_R0_data),
    .R0_en(mem_0_235_R0_en)
  );
  split_mem_0_ext mem_0_236 (
    .W0_addr(mem_0_236_W0_addr),
    .W0_clk(mem_0_236_W0_clk),
    .W0_data(mem_0_236_W0_data),
    .W0_en(mem_0_236_W0_en),
    .W0_mask(mem_0_236_W0_mask),
    .R0_addr(mem_0_236_R0_addr),
    .R0_clk(mem_0_236_R0_clk),
    .R0_data(mem_0_236_R0_data),
    .R0_en(mem_0_236_R0_en)
  );
  split_mem_0_ext mem_0_237 (
    .W0_addr(mem_0_237_W0_addr),
    .W0_clk(mem_0_237_W0_clk),
    .W0_data(mem_0_237_W0_data),
    .W0_en(mem_0_237_W0_en),
    .W0_mask(mem_0_237_W0_mask),
    .R0_addr(mem_0_237_R0_addr),
    .R0_clk(mem_0_237_R0_clk),
    .R0_data(mem_0_237_R0_data),
    .R0_en(mem_0_237_R0_en)
  );
  split_mem_0_ext mem_0_238 (
    .W0_addr(mem_0_238_W0_addr),
    .W0_clk(mem_0_238_W0_clk),
    .W0_data(mem_0_238_W0_data),
    .W0_en(mem_0_238_W0_en),
    .W0_mask(mem_0_238_W0_mask),
    .R0_addr(mem_0_238_R0_addr),
    .R0_clk(mem_0_238_R0_clk),
    .R0_data(mem_0_238_R0_data),
    .R0_en(mem_0_238_R0_en)
  );
  split_mem_0_ext mem_0_239 (
    .W0_addr(mem_0_239_W0_addr),
    .W0_clk(mem_0_239_W0_clk),
    .W0_data(mem_0_239_W0_data),
    .W0_en(mem_0_239_W0_en),
    .W0_mask(mem_0_239_W0_mask),
    .R0_addr(mem_0_239_R0_addr),
    .R0_clk(mem_0_239_R0_clk),
    .R0_data(mem_0_239_R0_data),
    .R0_en(mem_0_239_R0_en)
  );
  split_mem_0_ext mem_0_240 (
    .W0_addr(mem_0_240_W0_addr),
    .W0_clk(mem_0_240_W0_clk),
    .W0_data(mem_0_240_W0_data),
    .W0_en(mem_0_240_W0_en),
    .W0_mask(mem_0_240_W0_mask),
    .R0_addr(mem_0_240_R0_addr),
    .R0_clk(mem_0_240_R0_clk),
    .R0_data(mem_0_240_R0_data),
    .R0_en(mem_0_240_R0_en)
  );
  split_mem_0_ext mem_0_241 (
    .W0_addr(mem_0_241_W0_addr),
    .W0_clk(mem_0_241_W0_clk),
    .W0_data(mem_0_241_W0_data),
    .W0_en(mem_0_241_W0_en),
    .W0_mask(mem_0_241_W0_mask),
    .R0_addr(mem_0_241_R0_addr),
    .R0_clk(mem_0_241_R0_clk),
    .R0_data(mem_0_241_R0_data),
    .R0_en(mem_0_241_R0_en)
  );
  split_mem_0_ext mem_0_242 (
    .W0_addr(mem_0_242_W0_addr),
    .W0_clk(mem_0_242_W0_clk),
    .W0_data(mem_0_242_W0_data),
    .W0_en(mem_0_242_W0_en),
    .W0_mask(mem_0_242_W0_mask),
    .R0_addr(mem_0_242_R0_addr),
    .R0_clk(mem_0_242_R0_clk),
    .R0_data(mem_0_242_R0_data),
    .R0_en(mem_0_242_R0_en)
  );
  split_mem_0_ext mem_0_243 (
    .W0_addr(mem_0_243_W0_addr),
    .W0_clk(mem_0_243_W0_clk),
    .W0_data(mem_0_243_W0_data),
    .W0_en(mem_0_243_W0_en),
    .W0_mask(mem_0_243_W0_mask),
    .R0_addr(mem_0_243_R0_addr),
    .R0_clk(mem_0_243_R0_clk),
    .R0_data(mem_0_243_R0_data),
    .R0_en(mem_0_243_R0_en)
  );
  split_mem_0_ext mem_0_244 (
    .W0_addr(mem_0_244_W0_addr),
    .W0_clk(mem_0_244_W0_clk),
    .W0_data(mem_0_244_W0_data),
    .W0_en(mem_0_244_W0_en),
    .W0_mask(mem_0_244_W0_mask),
    .R0_addr(mem_0_244_R0_addr),
    .R0_clk(mem_0_244_R0_clk),
    .R0_data(mem_0_244_R0_data),
    .R0_en(mem_0_244_R0_en)
  );
  split_mem_0_ext mem_0_245 (
    .W0_addr(mem_0_245_W0_addr),
    .W0_clk(mem_0_245_W0_clk),
    .W0_data(mem_0_245_W0_data),
    .W0_en(mem_0_245_W0_en),
    .W0_mask(mem_0_245_W0_mask),
    .R0_addr(mem_0_245_R0_addr),
    .R0_clk(mem_0_245_R0_clk),
    .R0_data(mem_0_245_R0_data),
    .R0_en(mem_0_245_R0_en)
  );
  split_mem_0_ext mem_0_246 (
    .W0_addr(mem_0_246_W0_addr),
    .W0_clk(mem_0_246_W0_clk),
    .W0_data(mem_0_246_W0_data),
    .W0_en(mem_0_246_W0_en),
    .W0_mask(mem_0_246_W0_mask),
    .R0_addr(mem_0_246_R0_addr),
    .R0_clk(mem_0_246_R0_clk),
    .R0_data(mem_0_246_R0_data),
    .R0_en(mem_0_246_R0_en)
  );
  split_mem_0_ext mem_0_247 (
    .W0_addr(mem_0_247_W0_addr),
    .W0_clk(mem_0_247_W0_clk),
    .W0_data(mem_0_247_W0_data),
    .W0_en(mem_0_247_W0_en),
    .W0_mask(mem_0_247_W0_mask),
    .R0_addr(mem_0_247_R0_addr),
    .R0_clk(mem_0_247_R0_clk),
    .R0_data(mem_0_247_R0_data),
    .R0_en(mem_0_247_R0_en)
  );
  split_mem_0_ext mem_0_248 (
    .W0_addr(mem_0_248_W0_addr),
    .W0_clk(mem_0_248_W0_clk),
    .W0_data(mem_0_248_W0_data),
    .W0_en(mem_0_248_W0_en),
    .W0_mask(mem_0_248_W0_mask),
    .R0_addr(mem_0_248_R0_addr),
    .R0_clk(mem_0_248_R0_clk),
    .R0_data(mem_0_248_R0_data),
    .R0_en(mem_0_248_R0_en)
  );
  split_mem_0_ext mem_0_249 (
    .W0_addr(mem_0_249_W0_addr),
    .W0_clk(mem_0_249_W0_clk),
    .W0_data(mem_0_249_W0_data),
    .W0_en(mem_0_249_W0_en),
    .W0_mask(mem_0_249_W0_mask),
    .R0_addr(mem_0_249_R0_addr),
    .R0_clk(mem_0_249_R0_clk),
    .R0_data(mem_0_249_R0_data),
    .R0_en(mem_0_249_R0_en)
  );
  split_mem_0_ext mem_0_250 (
    .W0_addr(mem_0_250_W0_addr),
    .W0_clk(mem_0_250_W0_clk),
    .W0_data(mem_0_250_W0_data),
    .W0_en(mem_0_250_W0_en),
    .W0_mask(mem_0_250_W0_mask),
    .R0_addr(mem_0_250_R0_addr),
    .R0_clk(mem_0_250_R0_clk),
    .R0_data(mem_0_250_R0_data),
    .R0_en(mem_0_250_R0_en)
  );
  split_mem_0_ext mem_0_251 (
    .W0_addr(mem_0_251_W0_addr),
    .W0_clk(mem_0_251_W0_clk),
    .W0_data(mem_0_251_W0_data),
    .W0_en(mem_0_251_W0_en),
    .W0_mask(mem_0_251_W0_mask),
    .R0_addr(mem_0_251_R0_addr),
    .R0_clk(mem_0_251_R0_clk),
    .R0_data(mem_0_251_R0_data),
    .R0_en(mem_0_251_R0_en)
  );
  split_mem_0_ext mem_0_252 (
    .W0_addr(mem_0_252_W0_addr),
    .W0_clk(mem_0_252_W0_clk),
    .W0_data(mem_0_252_W0_data),
    .W0_en(mem_0_252_W0_en),
    .W0_mask(mem_0_252_W0_mask),
    .R0_addr(mem_0_252_R0_addr),
    .R0_clk(mem_0_252_R0_clk),
    .R0_data(mem_0_252_R0_data),
    .R0_en(mem_0_252_R0_en)
  );
  split_mem_0_ext mem_0_253 (
    .W0_addr(mem_0_253_W0_addr),
    .W0_clk(mem_0_253_W0_clk),
    .W0_data(mem_0_253_W0_data),
    .W0_en(mem_0_253_W0_en),
    .W0_mask(mem_0_253_W0_mask),
    .R0_addr(mem_0_253_R0_addr),
    .R0_clk(mem_0_253_R0_clk),
    .R0_data(mem_0_253_R0_data),
    .R0_en(mem_0_253_R0_en)
  );
  split_mem_0_ext mem_0_254 (
    .W0_addr(mem_0_254_W0_addr),
    .W0_clk(mem_0_254_W0_clk),
    .W0_data(mem_0_254_W0_data),
    .W0_en(mem_0_254_W0_en),
    .W0_mask(mem_0_254_W0_mask),
    .R0_addr(mem_0_254_R0_addr),
    .R0_clk(mem_0_254_R0_clk),
    .R0_data(mem_0_254_R0_data),
    .R0_en(mem_0_254_R0_en)
  );
  split_mem_0_ext mem_0_255 (
    .W0_addr(mem_0_255_W0_addr),
    .W0_clk(mem_0_255_W0_clk),
    .W0_data(mem_0_255_W0_data),
    .W0_en(mem_0_255_W0_en),
    .W0_mask(mem_0_255_W0_mask),
    .R0_addr(mem_0_255_R0_addr),
    .R0_clk(mem_0_255_R0_clk),
    .R0_data(mem_0_255_R0_data),
    .R0_en(mem_0_255_R0_en)
  );
  assign R0_data = {R0_data_0_255,_GEN_253};
  assign mem_0_0_W0_addr = W0_addr;
  assign mem_0_0_W0_clk = W0_clk;
  assign mem_0_0_W0_data = W0_data[7:0];
  assign mem_0_0_W0_en = W0_en;
  assign mem_0_0_W0_mask = W0_mask[0];
  assign mem_0_0_R0_addr = R0_addr;
  assign mem_0_0_R0_clk = R0_clk;
  assign mem_0_0_R0_en = R0_en;
  assign mem_0_1_W0_addr = W0_addr;
  assign mem_0_1_W0_clk = W0_clk;
  assign mem_0_1_W0_data = W0_data[15:8];
  assign mem_0_1_W0_en = W0_en;
  assign mem_0_1_W0_mask = W0_mask[1];
  assign mem_0_1_R0_addr = R0_addr;
  assign mem_0_1_R0_clk = R0_clk;
  assign mem_0_1_R0_en = R0_en;
  assign mem_0_2_W0_addr = W0_addr;
  assign mem_0_2_W0_clk = W0_clk;
  assign mem_0_2_W0_data = W0_data[23:16];
  assign mem_0_2_W0_en = W0_en;
  assign mem_0_2_W0_mask = W0_mask[2];
  assign mem_0_2_R0_addr = R0_addr;
  assign mem_0_2_R0_clk = R0_clk;
  assign mem_0_2_R0_en = R0_en;
  assign mem_0_3_W0_addr = W0_addr;
  assign mem_0_3_W0_clk = W0_clk;
  assign mem_0_3_W0_data = W0_data[31:24];
  assign mem_0_3_W0_en = W0_en;
  assign mem_0_3_W0_mask = W0_mask[3];
  assign mem_0_3_R0_addr = R0_addr;
  assign mem_0_3_R0_clk = R0_clk;
  assign mem_0_3_R0_en = R0_en;
  assign mem_0_4_W0_addr = W0_addr;
  assign mem_0_4_W0_clk = W0_clk;
  assign mem_0_4_W0_data = W0_data[39:32];
  assign mem_0_4_W0_en = W0_en;
  assign mem_0_4_W0_mask = W0_mask[4];
  assign mem_0_4_R0_addr = R0_addr;
  assign mem_0_4_R0_clk = R0_clk;
  assign mem_0_4_R0_en = R0_en;
  assign mem_0_5_W0_addr = W0_addr;
  assign mem_0_5_W0_clk = W0_clk;
  assign mem_0_5_W0_data = W0_data[47:40];
  assign mem_0_5_W0_en = W0_en;
  assign mem_0_5_W0_mask = W0_mask[5];
  assign mem_0_5_R0_addr = R0_addr;
  assign mem_0_5_R0_clk = R0_clk;
  assign mem_0_5_R0_en = R0_en;
  assign mem_0_6_W0_addr = W0_addr;
  assign mem_0_6_W0_clk = W0_clk;
  assign mem_0_6_W0_data = W0_data[55:48];
  assign mem_0_6_W0_en = W0_en;
  assign mem_0_6_W0_mask = W0_mask[6];
  assign mem_0_6_R0_addr = R0_addr;
  assign mem_0_6_R0_clk = R0_clk;
  assign mem_0_6_R0_en = R0_en;
  assign mem_0_7_W0_addr = W0_addr;
  assign mem_0_7_W0_clk = W0_clk;
  assign mem_0_7_W0_data = W0_data[63:56];
  assign mem_0_7_W0_en = W0_en;
  assign mem_0_7_W0_mask = W0_mask[7];
  assign mem_0_7_R0_addr = R0_addr;
  assign mem_0_7_R0_clk = R0_clk;
  assign mem_0_7_R0_en = R0_en;
  assign mem_0_8_W0_addr = W0_addr;
  assign mem_0_8_W0_clk = W0_clk;
  assign mem_0_8_W0_data = W0_data[71:64];
  assign mem_0_8_W0_en = W0_en;
  assign mem_0_8_W0_mask = W0_mask[8];
  assign mem_0_8_R0_addr = R0_addr;
  assign mem_0_8_R0_clk = R0_clk;
  assign mem_0_8_R0_en = R0_en;
  assign mem_0_9_W0_addr = W0_addr;
  assign mem_0_9_W0_clk = W0_clk;
  assign mem_0_9_W0_data = W0_data[79:72];
  assign mem_0_9_W0_en = W0_en;
  assign mem_0_9_W0_mask = W0_mask[9];
  assign mem_0_9_R0_addr = R0_addr;
  assign mem_0_9_R0_clk = R0_clk;
  assign mem_0_9_R0_en = R0_en;
  assign mem_0_10_W0_addr = W0_addr;
  assign mem_0_10_W0_clk = W0_clk;
  assign mem_0_10_W0_data = W0_data[87:80];
  assign mem_0_10_W0_en = W0_en;
  assign mem_0_10_W0_mask = W0_mask[10];
  assign mem_0_10_R0_addr = R0_addr;
  assign mem_0_10_R0_clk = R0_clk;
  assign mem_0_10_R0_en = R0_en;
  assign mem_0_11_W0_addr = W0_addr;
  assign mem_0_11_W0_clk = W0_clk;
  assign mem_0_11_W0_data = W0_data[95:88];
  assign mem_0_11_W0_en = W0_en;
  assign mem_0_11_W0_mask = W0_mask[11];
  assign mem_0_11_R0_addr = R0_addr;
  assign mem_0_11_R0_clk = R0_clk;
  assign mem_0_11_R0_en = R0_en;
  assign mem_0_12_W0_addr = W0_addr;
  assign mem_0_12_W0_clk = W0_clk;
  assign mem_0_12_W0_data = W0_data[103:96];
  assign mem_0_12_W0_en = W0_en;
  assign mem_0_12_W0_mask = W0_mask[12];
  assign mem_0_12_R0_addr = R0_addr;
  assign mem_0_12_R0_clk = R0_clk;
  assign mem_0_12_R0_en = R0_en;
  assign mem_0_13_W0_addr = W0_addr;
  assign mem_0_13_W0_clk = W0_clk;
  assign mem_0_13_W0_data = W0_data[111:104];
  assign mem_0_13_W0_en = W0_en;
  assign mem_0_13_W0_mask = W0_mask[13];
  assign mem_0_13_R0_addr = R0_addr;
  assign mem_0_13_R0_clk = R0_clk;
  assign mem_0_13_R0_en = R0_en;
  assign mem_0_14_W0_addr = W0_addr;
  assign mem_0_14_W0_clk = W0_clk;
  assign mem_0_14_W0_data = W0_data[119:112];
  assign mem_0_14_W0_en = W0_en;
  assign mem_0_14_W0_mask = W0_mask[14];
  assign mem_0_14_R0_addr = R0_addr;
  assign mem_0_14_R0_clk = R0_clk;
  assign mem_0_14_R0_en = R0_en;
  assign mem_0_15_W0_addr = W0_addr;
  assign mem_0_15_W0_clk = W0_clk;
  assign mem_0_15_W0_data = W0_data[127:120];
  assign mem_0_15_W0_en = W0_en;
  assign mem_0_15_W0_mask = W0_mask[15];
  assign mem_0_15_R0_addr = R0_addr;
  assign mem_0_15_R0_clk = R0_clk;
  assign mem_0_15_R0_en = R0_en;
  assign mem_0_16_W0_addr = W0_addr;
  assign mem_0_16_W0_clk = W0_clk;
  assign mem_0_16_W0_data = W0_data[135:128];
  assign mem_0_16_W0_en = W0_en;
  assign mem_0_16_W0_mask = W0_mask[16];
  assign mem_0_16_R0_addr = R0_addr;
  assign mem_0_16_R0_clk = R0_clk;
  assign mem_0_16_R0_en = R0_en;
  assign mem_0_17_W0_addr = W0_addr;
  assign mem_0_17_W0_clk = W0_clk;
  assign mem_0_17_W0_data = W0_data[143:136];
  assign mem_0_17_W0_en = W0_en;
  assign mem_0_17_W0_mask = W0_mask[17];
  assign mem_0_17_R0_addr = R0_addr;
  assign mem_0_17_R0_clk = R0_clk;
  assign mem_0_17_R0_en = R0_en;
  assign mem_0_18_W0_addr = W0_addr;
  assign mem_0_18_W0_clk = W0_clk;
  assign mem_0_18_W0_data = W0_data[151:144];
  assign mem_0_18_W0_en = W0_en;
  assign mem_0_18_W0_mask = W0_mask[18];
  assign mem_0_18_R0_addr = R0_addr;
  assign mem_0_18_R0_clk = R0_clk;
  assign mem_0_18_R0_en = R0_en;
  assign mem_0_19_W0_addr = W0_addr;
  assign mem_0_19_W0_clk = W0_clk;
  assign mem_0_19_W0_data = W0_data[159:152];
  assign mem_0_19_W0_en = W0_en;
  assign mem_0_19_W0_mask = W0_mask[19];
  assign mem_0_19_R0_addr = R0_addr;
  assign mem_0_19_R0_clk = R0_clk;
  assign mem_0_19_R0_en = R0_en;
  assign mem_0_20_W0_addr = W0_addr;
  assign mem_0_20_W0_clk = W0_clk;
  assign mem_0_20_W0_data = W0_data[167:160];
  assign mem_0_20_W0_en = W0_en;
  assign mem_0_20_W0_mask = W0_mask[20];
  assign mem_0_20_R0_addr = R0_addr;
  assign mem_0_20_R0_clk = R0_clk;
  assign mem_0_20_R0_en = R0_en;
  assign mem_0_21_W0_addr = W0_addr;
  assign mem_0_21_W0_clk = W0_clk;
  assign mem_0_21_W0_data = W0_data[175:168];
  assign mem_0_21_W0_en = W0_en;
  assign mem_0_21_W0_mask = W0_mask[21];
  assign mem_0_21_R0_addr = R0_addr;
  assign mem_0_21_R0_clk = R0_clk;
  assign mem_0_21_R0_en = R0_en;
  assign mem_0_22_W0_addr = W0_addr;
  assign mem_0_22_W0_clk = W0_clk;
  assign mem_0_22_W0_data = W0_data[183:176];
  assign mem_0_22_W0_en = W0_en;
  assign mem_0_22_W0_mask = W0_mask[22];
  assign mem_0_22_R0_addr = R0_addr;
  assign mem_0_22_R0_clk = R0_clk;
  assign mem_0_22_R0_en = R0_en;
  assign mem_0_23_W0_addr = W0_addr;
  assign mem_0_23_W0_clk = W0_clk;
  assign mem_0_23_W0_data = W0_data[191:184];
  assign mem_0_23_W0_en = W0_en;
  assign mem_0_23_W0_mask = W0_mask[23];
  assign mem_0_23_R0_addr = R0_addr;
  assign mem_0_23_R0_clk = R0_clk;
  assign mem_0_23_R0_en = R0_en;
  assign mem_0_24_W0_addr = W0_addr;
  assign mem_0_24_W0_clk = W0_clk;
  assign mem_0_24_W0_data = W0_data[199:192];
  assign mem_0_24_W0_en = W0_en;
  assign mem_0_24_W0_mask = W0_mask[24];
  assign mem_0_24_R0_addr = R0_addr;
  assign mem_0_24_R0_clk = R0_clk;
  assign mem_0_24_R0_en = R0_en;
  assign mem_0_25_W0_addr = W0_addr;
  assign mem_0_25_W0_clk = W0_clk;
  assign mem_0_25_W0_data = W0_data[207:200];
  assign mem_0_25_W0_en = W0_en;
  assign mem_0_25_W0_mask = W0_mask[25];
  assign mem_0_25_R0_addr = R0_addr;
  assign mem_0_25_R0_clk = R0_clk;
  assign mem_0_25_R0_en = R0_en;
  assign mem_0_26_W0_addr = W0_addr;
  assign mem_0_26_W0_clk = W0_clk;
  assign mem_0_26_W0_data = W0_data[215:208];
  assign mem_0_26_W0_en = W0_en;
  assign mem_0_26_W0_mask = W0_mask[26];
  assign mem_0_26_R0_addr = R0_addr;
  assign mem_0_26_R0_clk = R0_clk;
  assign mem_0_26_R0_en = R0_en;
  assign mem_0_27_W0_addr = W0_addr;
  assign mem_0_27_W0_clk = W0_clk;
  assign mem_0_27_W0_data = W0_data[223:216];
  assign mem_0_27_W0_en = W0_en;
  assign mem_0_27_W0_mask = W0_mask[27];
  assign mem_0_27_R0_addr = R0_addr;
  assign mem_0_27_R0_clk = R0_clk;
  assign mem_0_27_R0_en = R0_en;
  assign mem_0_28_W0_addr = W0_addr;
  assign mem_0_28_W0_clk = W0_clk;
  assign mem_0_28_W0_data = W0_data[231:224];
  assign mem_0_28_W0_en = W0_en;
  assign mem_0_28_W0_mask = W0_mask[28];
  assign mem_0_28_R0_addr = R0_addr;
  assign mem_0_28_R0_clk = R0_clk;
  assign mem_0_28_R0_en = R0_en;
  assign mem_0_29_W0_addr = W0_addr;
  assign mem_0_29_W0_clk = W0_clk;
  assign mem_0_29_W0_data = W0_data[239:232];
  assign mem_0_29_W0_en = W0_en;
  assign mem_0_29_W0_mask = W0_mask[29];
  assign mem_0_29_R0_addr = R0_addr;
  assign mem_0_29_R0_clk = R0_clk;
  assign mem_0_29_R0_en = R0_en;
  assign mem_0_30_W0_addr = W0_addr;
  assign mem_0_30_W0_clk = W0_clk;
  assign mem_0_30_W0_data = W0_data[247:240];
  assign mem_0_30_W0_en = W0_en;
  assign mem_0_30_W0_mask = W0_mask[30];
  assign mem_0_30_R0_addr = R0_addr;
  assign mem_0_30_R0_clk = R0_clk;
  assign mem_0_30_R0_en = R0_en;
  assign mem_0_31_W0_addr = W0_addr;
  assign mem_0_31_W0_clk = W0_clk;
  assign mem_0_31_W0_data = W0_data[255:248];
  assign mem_0_31_W0_en = W0_en;
  assign mem_0_31_W0_mask = W0_mask[31];
  assign mem_0_31_R0_addr = R0_addr;
  assign mem_0_31_R0_clk = R0_clk;
  assign mem_0_31_R0_en = R0_en;
  assign mem_0_32_W0_addr = W0_addr;
  assign mem_0_32_W0_clk = W0_clk;
  assign mem_0_32_W0_data = W0_data[263:256];
  assign mem_0_32_W0_en = W0_en;
  assign mem_0_32_W0_mask = W0_mask[32];
  assign mem_0_32_R0_addr = R0_addr;
  assign mem_0_32_R0_clk = R0_clk;
  assign mem_0_32_R0_en = R0_en;
  assign mem_0_33_W0_addr = W0_addr;
  assign mem_0_33_W0_clk = W0_clk;
  assign mem_0_33_W0_data = W0_data[271:264];
  assign mem_0_33_W0_en = W0_en;
  assign mem_0_33_W0_mask = W0_mask[33];
  assign mem_0_33_R0_addr = R0_addr;
  assign mem_0_33_R0_clk = R0_clk;
  assign mem_0_33_R0_en = R0_en;
  assign mem_0_34_W0_addr = W0_addr;
  assign mem_0_34_W0_clk = W0_clk;
  assign mem_0_34_W0_data = W0_data[279:272];
  assign mem_0_34_W0_en = W0_en;
  assign mem_0_34_W0_mask = W0_mask[34];
  assign mem_0_34_R0_addr = R0_addr;
  assign mem_0_34_R0_clk = R0_clk;
  assign mem_0_34_R0_en = R0_en;
  assign mem_0_35_W0_addr = W0_addr;
  assign mem_0_35_W0_clk = W0_clk;
  assign mem_0_35_W0_data = W0_data[287:280];
  assign mem_0_35_W0_en = W0_en;
  assign mem_0_35_W0_mask = W0_mask[35];
  assign mem_0_35_R0_addr = R0_addr;
  assign mem_0_35_R0_clk = R0_clk;
  assign mem_0_35_R0_en = R0_en;
  assign mem_0_36_W0_addr = W0_addr;
  assign mem_0_36_W0_clk = W0_clk;
  assign mem_0_36_W0_data = W0_data[295:288];
  assign mem_0_36_W0_en = W0_en;
  assign mem_0_36_W0_mask = W0_mask[36];
  assign mem_0_36_R0_addr = R0_addr;
  assign mem_0_36_R0_clk = R0_clk;
  assign mem_0_36_R0_en = R0_en;
  assign mem_0_37_W0_addr = W0_addr;
  assign mem_0_37_W0_clk = W0_clk;
  assign mem_0_37_W0_data = W0_data[303:296];
  assign mem_0_37_W0_en = W0_en;
  assign mem_0_37_W0_mask = W0_mask[37];
  assign mem_0_37_R0_addr = R0_addr;
  assign mem_0_37_R0_clk = R0_clk;
  assign mem_0_37_R0_en = R0_en;
  assign mem_0_38_W0_addr = W0_addr;
  assign mem_0_38_W0_clk = W0_clk;
  assign mem_0_38_W0_data = W0_data[311:304];
  assign mem_0_38_W0_en = W0_en;
  assign mem_0_38_W0_mask = W0_mask[38];
  assign mem_0_38_R0_addr = R0_addr;
  assign mem_0_38_R0_clk = R0_clk;
  assign mem_0_38_R0_en = R0_en;
  assign mem_0_39_W0_addr = W0_addr;
  assign mem_0_39_W0_clk = W0_clk;
  assign mem_0_39_W0_data = W0_data[319:312];
  assign mem_0_39_W0_en = W0_en;
  assign mem_0_39_W0_mask = W0_mask[39];
  assign mem_0_39_R0_addr = R0_addr;
  assign mem_0_39_R0_clk = R0_clk;
  assign mem_0_39_R0_en = R0_en;
  assign mem_0_40_W0_addr = W0_addr;
  assign mem_0_40_W0_clk = W0_clk;
  assign mem_0_40_W0_data = W0_data[327:320];
  assign mem_0_40_W0_en = W0_en;
  assign mem_0_40_W0_mask = W0_mask[40];
  assign mem_0_40_R0_addr = R0_addr;
  assign mem_0_40_R0_clk = R0_clk;
  assign mem_0_40_R0_en = R0_en;
  assign mem_0_41_W0_addr = W0_addr;
  assign mem_0_41_W0_clk = W0_clk;
  assign mem_0_41_W0_data = W0_data[335:328];
  assign mem_0_41_W0_en = W0_en;
  assign mem_0_41_W0_mask = W0_mask[41];
  assign mem_0_41_R0_addr = R0_addr;
  assign mem_0_41_R0_clk = R0_clk;
  assign mem_0_41_R0_en = R0_en;
  assign mem_0_42_W0_addr = W0_addr;
  assign mem_0_42_W0_clk = W0_clk;
  assign mem_0_42_W0_data = W0_data[343:336];
  assign mem_0_42_W0_en = W0_en;
  assign mem_0_42_W0_mask = W0_mask[42];
  assign mem_0_42_R0_addr = R0_addr;
  assign mem_0_42_R0_clk = R0_clk;
  assign mem_0_42_R0_en = R0_en;
  assign mem_0_43_W0_addr = W0_addr;
  assign mem_0_43_W0_clk = W0_clk;
  assign mem_0_43_W0_data = W0_data[351:344];
  assign mem_0_43_W0_en = W0_en;
  assign mem_0_43_W0_mask = W0_mask[43];
  assign mem_0_43_R0_addr = R0_addr;
  assign mem_0_43_R0_clk = R0_clk;
  assign mem_0_43_R0_en = R0_en;
  assign mem_0_44_W0_addr = W0_addr;
  assign mem_0_44_W0_clk = W0_clk;
  assign mem_0_44_W0_data = W0_data[359:352];
  assign mem_0_44_W0_en = W0_en;
  assign mem_0_44_W0_mask = W0_mask[44];
  assign mem_0_44_R0_addr = R0_addr;
  assign mem_0_44_R0_clk = R0_clk;
  assign mem_0_44_R0_en = R0_en;
  assign mem_0_45_W0_addr = W0_addr;
  assign mem_0_45_W0_clk = W0_clk;
  assign mem_0_45_W0_data = W0_data[367:360];
  assign mem_0_45_W0_en = W0_en;
  assign mem_0_45_W0_mask = W0_mask[45];
  assign mem_0_45_R0_addr = R0_addr;
  assign mem_0_45_R0_clk = R0_clk;
  assign mem_0_45_R0_en = R0_en;
  assign mem_0_46_W0_addr = W0_addr;
  assign mem_0_46_W0_clk = W0_clk;
  assign mem_0_46_W0_data = W0_data[375:368];
  assign mem_0_46_W0_en = W0_en;
  assign mem_0_46_W0_mask = W0_mask[46];
  assign mem_0_46_R0_addr = R0_addr;
  assign mem_0_46_R0_clk = R0_clk;
  assign mem_0_46_R0_en = R0_en;
  assign mem_0_47_W0_addr = W0_addr;
  assign mem_0_47_W0_clk = W0_clk;
  assign mem_0_47_W0_data = W0_data[383:376];
  assign mem_0_47_W0_en = W0_en;
  assign mem_0_47_W0_mask = W0_mask[47];
  assign mem_0_47_R0_addr = R0_addr;
  assign mem_0_47_R0_clk = R0_clk;
  assign mem_0_47_R0_en = R0_en;
  assign mem_0_48_W0_addr = W0_addr;
  assign mem_0_48_W0_clk = W0_clk;
  assign mem_0_48_W0_data = W0_data[391:384];
  assign mem_0_48_W0_en = W0_en;
  assign mem_0_48_W0_mask = W0_mask[48];
  assign mem_0_48_R0_addr = R0_addr;
  assign mem_0_48_R0_clk = R0_clk;
  assign mem_0_48_R0_en = R0_en;
  assign mem_0_49_W0_addr = W0_addr;
  assign mem_0_49_W0_clk = W0_clk;
  assign mem_0_49_W0_data = W0_data[399:392];
  assign mem_0_49_W0_en = W0_en;
  assign mem_0_49_W0_mask = W0_mask[49];
  assign mem_0_49_R0_addr = R0_addr;
  assign mem_0_49_R0_clk = R0_clk;
  assign mem_0_49_R0_en = R0_en;
  assign mem_0_50_W0_addr = W0_addr;
  assign mem_0_50_W0_clk = W0_clk;
  assign mem_0_50_W0_data = W0_data[407:400];
  assign mem_0_50_W0_en = W0_en;
  assign mem_0_50_W0_mask = W0_mask[50];
  assign mem_0_50_R0_addr = R0_addr;
  assign mem_0_50_R0_clk = R0_clk;
  assign mem_0_50_R0_en = R0_en;
  assign mem_0_51_W0_addr = W0_addr;
  assign mem_0_51_W0_clk = W0_clk;
  assign mem_0_51_W0_data = W0_data[415:408];
  assign mem_0_51_W0_en = W0_en;
  assign mem_0_51_W0_mask = W0_mask[51];
  assign mem_0_51_R0_addr = R0_addr;
  assign mem_0_51_R0_clk = R0_clk;
  assign mem_0_51_R0_en = R0_en;
  assign mem_0_52_W0_addr = W0_addr;
  assign mem_0_52_W0_clk = W0_clk;
  assign mem_0_52_W0_data = W0_data[423:416];
  assign mem_0_52_W0_en = W0_en;
  assign mem_0_52_W0_mask = W0_mask[52];
  assign mem_0_52_R0_addr = R0_addr;
  assign mem_0_52_R0_clk = R0_clk;
  assign mem_0_52_R0_en = R0_en;
  assign mem_0_53_W0_addr = W0_addr;
  assign mem_0_53_W0_clk = W0_clk;
  assign mem_0_53_W0_data = W0_data[431:424];
  assign mem_0_53_W0_en = W0_en;
  assign mem_0_53_W0_mask = W0_mask[53];
  assign mem_0_53_R0_addr = R0_addr;
  assign mem_0_53_R0_clk = R0_clk;
  assign mem_0_53_R0_en = R0_en;
  assign mem_0_54_W0_addr = W0_addr;
  assign mem_0_54_W0_clk = W0_clk;
  assign mem_0_54_W0_data = W0_data[439:432];
  assign mem_0_54_W0_en = W0_en;
  assign mem_0_54_W0_mask = W0_mask[54];
  assign mem_0_54_R0_addr = R0_addr;
  assign mem_0_54_R0_clk = R0_clk;
  assign mem_0_54_R0_en = R0_en;
  assign mem_0_55_W0_addr = W0_addr;
  assign mem_0_55_W0_clk = W0_clk;
  assign mem_0_55_W0_data = W0_data[447:440];
  assign mem_0_55_W0_en = W0_en;
  assign mem_0_55_W0_mask = W0_mask[55];
  assign mem_0_55_R0_addr = R0_addr;
  assign mem_0_55_R0_clk = R0_clk;
  assign mem_0_55_R0_en = R0_en;
  assign mem_0_56_W0_addr = W0_addr;
  assign mem_0_56_W0_clk = W0_clk;
  assign mem_0_56_W0_data = W0_data[455:448];
  assign mem_0_56_W0_en = W0_en;
  assign mem_0_56_W0_mask = W0_mask[56];
  assign mem_0_56_R0_addr = R0_addr;
  assign mem_0_56_R0_clk = R0_clk;
  assign mem_0_56_R0_en = R0_en;
  assign mem_0_57_W0_addr = W0_addr;
  assign mem_0_57_W0_clk = W0_clk;
  assign mem_0_57_W0_data = W0_data[463:456];
  assign mem_0_57_W0_en = W0_en;
  assign mem_0_57_W0_mask = W0_mask[57];
  assign mem_0_57_R0_addr = R0_addr;
  assign mem_0_57_R0_clk = R0_clk;
  assign mem_0_57_R0_en = R0_en;
  assign mem_0_58_W0_addr = W0_addr;
  assign mem_0_58_W0_clk = W0_clk;
  assign mem_0_58_W0_data = W0_data[471:464];
  assign mem_0_58_W0_en = W0_en;
  assign mem_0_58_W0_mask = W0_mask[58];
  assign mem_0_58_R0_addr = R0_addr;
  assign mem_0_58_R0_clk = R0_clk;
  assign mem_0_58_R0_en = R0_en;
  assign mem_0_59_W0_addr = W0_addr;
  assign mem_0_59_W0_clk = W0_clk;
  assign mem_0_59_W0_data = W0_data[479:472];
  assign mem_0_59_W0_en = W0_en;
  assign mem_0_59_W0_mask = W0_mask[59];
  assign mem_0_59_R0_addr = R0_addr;
  assign mem_0_59_R0_clk = R0_clk;
  assign mem_0_59_R0_en = R0_en;
  assign mem_0_60_W0_addr = W0_addr;
  assign mem_0_60_W0_clk = W0_clk;
  assign mem_0_60_W0_data = W0_data[487:480];
  assign mem_0_60_W0_en = W0_en;
  assign mem_0_60_W0_mask = W0_mask[60];
  assign mem_0_60_R0_addr = R0_addr;
  assign mem_0_60_R0_clk = R0_clk;
  assign mem_0_60_R0_en = R0_en;
  assign mem_0_61_W0_addr = W0_addr;
  assign mem_0_61_W0_clk = W0_clk;
  assign mem_0_61_W0_data = W0_data[495:488];
  assign mem_0_61_W0_en = W0_en;
  assign mem_0_61_W0_mask = W0_mask[61];
  assign mem_0_61_R0_addr = R0_addr;
  assign mem_0_61_R0_clk = R0_clk;
  assign mem_0_61_R0_en = R0_en;
  assign mem_0_62_W0_addr = W0_addr;
  assign mem_0_62_W0_clk = W0_clk;
  assign mem_0_62_W0_data = W0_data[503:496];
  assign mem_0_62_W0_en = W0_en;
  assign mem_0_62_W0_mask = W0_mask[62];
  assign mem_0_62_R0_addr = R0_addr;
  assign mem_0_62_R0_clk = R0_clk;
  assign mem_0_62_R0_en = R0_en;
  assign mem_0_63_W0_addr = W0_addr;
  assign mem_0_63_W0_clk = W0_clk;
  assign mem_0_63_W0_data = W0_data[511:504];
  assign mem_0_63_W0_en = W0_en;
  assign mem_0_63_W0_mask = W0_mask[63];
  assign mem_0_63_R0_addr = R0_addr;
  assign mem_0_63_R0_clk = R0_clk;
  assign mem_0_63_R0_en = R0_en;
  assign mem_0_64_W0_addr = W0_addr;
  assign mem_0_64_W0_clk = W0_clk;
  assign mem_0_64_W0_data = W0_data[519:512];
  assign mem_0_64_W0_en = W0_en;
  assign mem_0_64_W0_mask = W0_mask[64];
  assign mem_0_64_R0_addr = R0_addr;
  assign mem_0_64_R0_clk = R0_clk;
  assign mem_0_64_R0_en = R0_en;
  assign mem_0_65_W0_addr = W0_addr;
  assign mem_0_65_W0_clk = W0_clk;
  assign mem_0_65_W0_data = W0_data[527:520];
  assign mem_0_65_W0_en = W0_en;
  assign mem_0_65_W0_mask = W0_mask[65];
  assign mem_0_65_R0_addr = R0_addr;
  assign mem_0_65_R0_clk = R0_clk;
  assign mem_0_65_R0_en = R0_en;
  assign mem_0_66_W0_addr = W0_addr;
  assign mem_0_66_W0_clk = W0_clk;
  assign mem_0_66_W0_data = W0_data[535:528];
  assign mem_0_66_W0_en = W0_en;
  assign mem_0_66_W0_mask = W0_mask[66];
  assign mem_0_66_R0_addr = R0_addr;
  assign mem_0_66_R0_clk = R0_clk;
  assign mem_0_66_R0_en = R0_en;
  assign mem_0_67_W0_addr = W0_addr;
  assign mem_0_67_W0_clk = W0_clk;
  assign mem_0_67_W0_data = W0_data[543:536];
  assign mem_0_67_W0_en = W0_en;
  assign mem_0_67_W0_mask = W0_mask[67];
  assign mem_0_67_R0_addr = R0_addr;
  assign mem_0_67_R0_clk = R0_clk;
  assign mem_0_67_R0_en = R0_en;
  assign mem_0_68_W0_addr = W0_addr;
  assign mem_0_68_W0_clk = W0_clk;
  assign mem_0_68_W0_data = W0_data[551:544];
  assign mem_0_68_W0_en = W0_en;
  assign mem_0_68_W0_mask = W0_mask[68];
  assign mem_0_68_R0_addr = R0_addr;
  assign mem_0_68_R0_clk = R0_clk;
  assign mem_0_68_R0_en = R0_en;
  assign mem_0_69_W0_addr = W0_addr;
  assign mem_0_69_W0_clk = W0_clk;
  assign mem_0_69_W0_data = W0_data[559:552];
  assign mem_0_69_W0_en = W0_en;
  assign mem_0_69_W0_mask = W0_mask[69];
  assign mem_0_69_R0_addr = R0_addr;
  assign mem_0_69_R0_clk = R0_clk;
  assign mem_0_69_R0_en = R0_en;
  assign mem_0_70_W0_addr = W0_addr;
  assign mem_0_70_W0_clk = W0_clk;
  assign mem_0_70_W0_data = W0_data[567:560];
  assign mem_0_70_W0_en = W0_en;
  assign mem_0_70_W0_mask = W0_mask[70];
  assign mem_0_70_R0_addr = R0_addr;
  assign mem_0_70_R0_clk = R0_clk;
  assign mem_0_70_R0_en = R0_en;
  assign mem_0_71_W0_addr = W0_addr;
  assign mem_0_71_W0_clk = W0_clk;
  assign mem_0_71_W0_data = W0_data[575:568];
  assign mem_0_71_W0_en = W0_en;
  assign mem_0_71_W0_mask = W0_mask[71];
  assign mem_0_71_R0_addr = R0_addr;
  assign mem_0_71_R0_clk = R0_clk;
  assign mem_0_71_R0_en = R0_en;
  assign mem_0_72_W0_addr = W0_addr;
  assign mem_0_72_W0_clk = W0_clk;
  assign mem_0_72_W0_data = W0_data[583:576];
  assign mem_0_72_W0_en = W0_en;
  assign mem_0_72_W0_mask = W0_mask[72];
  assign mem_0_72_R0_addr = R0_addr;
  assign mem_0_72_R0_clk = R0_clk;
  assign mem_0_72_R0_en = R0_en;
  assign mem_0_73_W0_addr = W0_addr;
  assign mem_0_73_W0_clk = W0_clk;
  assign mem_0_73_W0_data = W0_data[591:584];
  assign mem_0_73_W0_en = W0_en;
  assign mem_0_73_W0_mask = W0_mask[73];
  assign mem_0_73_R0_addr = R0_addr;
  assign mem_0_73_R0_clk = R0_clk;
  assign mem_0_73_R0_en = R0_en;
  assign mem_0_74_W0_addr = W0_addr;
  assign mem_0_74_W0_clk = W0_clk;
  assign mem_0_74_W0_data = W0_data[599:592];
  assign mem_0_74_W0_en = W0_en;
  assign mem_0_74_W0_mask = W0_mask[74];
  assign mem_0_74_R0_addr = R0_addr;
  assign mem_0_74_R0_clk = R0_clk;
  assign mem_0_74_R0_en = R0_en;
  assign mem_0_75_W0_addr = W0_addr;
  assign mem_0_75_W0_clk = W0_clk;
  assign mem_0_75_W0_data = W0_data[607:600];
  assign mem_0_75_W0_en = W0_en;
  assign mem_0_75_W0_mask = W0_mask[75];
  assign mem_0_75_R0_addr = R0_addr;
  assign mem_0_75_R0_clk = R0_clk;
  assign mem_0_75_R0_en = R0_en;
  assign mem_0_76_W0_addr = W0_addr;
  assign mem_0_76_W0_clk = W0_clk;
  assign mem_0_76_W0_data = W0_data[615:608];
  assign mem_0_76_W0_en = W0_en;
  assign mem_0_76_W0_mask = W0_mask[76];
  assign mem_0_76_R0_addr = R0_addr;
  assign mem_0_76_R0_clk = R0_clk;
  assign mem_0_76_R0_en = R0_en;
  assign mem_0_77_W0_addr = W0_addr;
  assign mem_0_77_W0_clk = W0_clk;
  assign mem_0_77_W0_data = W0_data[623:616];
  assign mem_0_77_W0_en = W0_en;
  assign mem_0_77_W0_mask = W0_mask[77];
  assign mem_0_77_R0_addr = R0_addr;
  assign mem_0_77_R0_clk = R0_clk;
  assign mem_0_77_R0_en = R0_en;
  assign mem_0_78_W0_addr = W0_addr;
  assign mem_0_78_W0_clk = W0_clk;
  assign mem_0_78_W0_data = W0_data[631:624];
  assign mem_0_78_W0_en = W0_en;
  assign mem_0_78_W0_mask = W0_mask[78];
  assign mem_0_78_R0_addr = R0_addr;
  assign mem_0_78_R0_clk = R0_clk;
  assign mem_0_78_R0_en = R0_en;
  assign mem_0_79_W0_addr = W0_addr;
  assign mem_0_79_W0_clk = W0_clk;
  assign mem_0_79_W0_data = W0_data[639:632];
  assign mem_0_79_W0_en = W0_en;
  assign mem_0_79_W0_mask = W0_mask[79];
  assign mem_0_79_R0_addr = R0_addr;
  assign mem_0_79_R0_clk = R0_clk;
  assign mem_0_79_R0_en = R0_en;
  assign mem_0_80_W0_addr = W0_addr;
  assign mem_0_80_W0_clk = W0_clk;
  assign mem_0_80_W0_data = W0_data[647:640];
  assign mem_0_80_W0_en = W0_en;
  assign mem_0_80_W0_mask = W0_mask[80];
  assign mem_0_80_R0_addr = R0_addr;
  assign mem_0_80_R0_clk = R0_clk;
  assign mem_0_80_R0_en = R0_en;
  assign mem_0_81_W0_addr = W0_addr;
  assign mem_0_81_W0_clk = W0_clk;
  assign mem_0_81_W0_data = W0_data[655:648];
  assign mem_0_81_W0_en = W0_en;
  assign mem_0_81_W0_mask = W0_mask[81];
  assign mem_0_81_R0_addr = R0_addr;
  assign mem_0_81_R0_clk = R0_clk;
  assign mem_0_81_R0_en = R0_en;
  assign mem_0_82_W0_addr = W0_addr;
  assign mem_0_82_W0_clk = W0_clk;
  assign mem_0_82_W0_data = W0_data[663:656];
  assign mem_0_82_W0_en = W0_en;
  assign mem_0_82_W0_mask = W0_mask[82];
  assign mem_0_82_R0_addr = R0_addr;
  assign mem_0_82_R0_clk = R0_clk;
  assign mem_0_82_R0_en = R0_en;
  assign mem_0_83_W0_addr = W0_addr;
  assign mem_0_83_W0_clk = W0_clk;
  assign mem_0_83_W0_data = W0_data[671:664];
  assign mem_0_83_W0_en = W0_en;
  assign mem_0_83_W0_mask = W0_mask[83];
  assign mem_0_83_R0_addr = R0_addr;
  assign mem_0_83_R0_clk = R0_clk;
  assign mem_0_83_R0_en = R0_en;
  assign mem_0_84_W0_addr = W0_addr;
  assign mem_0_84_W0_clk = W0_clk;
  assign mem_0_84_W0_data = W0_data[679:672];
  assign mem_0_84_W0_en = W0_en;
  assign mem_0_84_W0_mask = W0_mask[84];
  assign mem_0_84_R0_addr = R0_addr;
  assign mem_0_84_R0_clk = R0_clk;
  assign mem_0_84_R0_en = R0_en;
  assign mem_0_85_W0_addr = W0_addr;
  assign mem_0_85_W0_clk = W0_clk;
  assign mem_0_85_W0_data = W0_data[687:680];
  assign mem_0_85_W0_en = W0_en;
  assign mem_0_85_W0_mask = W0_mask[85];
  assign mem_0_85_R0_addr = R0_addr;
  assign mem_0_85_R0_clk = R0_clk;
  assign mem_0_85_R0_en = R0_en;
  assign mem_0_86_W0_addr = W0_addr;
  assign mem_0_86_W0_clk = W0_clk;
  assign mem_0_86_W0_data = W0_data[695:688];
  assign mem_0_86_W0_en = W0_en;
  assign mem_0_86_W0_mask = W0_mask[86];
  assign mem_0_86_R0_addr = R0_addr;
  assign mem_0_86_R0_clk = R0_clk;
  assign mem_0_86_R0_en = R0_en;
  assign mem_0_87_W0_addr = W0_addr;
  assign mem_0_87_W0_clk = W0_clk;
  assign mem_0_87_W0_data = W0_data[703:696];
  assign mem_0_87_W0_en = W0_en;
  assign mem_0_87_W0_mask = W0_mask[87];
  assign mem_0_87_R0_addr = R0_addr;
  assign mem_0_87_R0_clk = R0_clk;
  assign mem_0_87_R0_en = R0_en;
  assign mem_0_88_W0_addr = W0_addr;
  assign mem_0_88_W0_clk = W0_clk;
  assign mem_0_88_W0_data = W0_data[711:704];
  assign mem_0_88_W0_en = W0_en;
  assign mem_0_88_W0_mask = W0_mask[88];
  assign mem_0_88_R0_addr = R0_addr;
  assign mem_0_88_R0_clk = R0_clk;
  assign mem_0_88_R0_en = R0_en;
  assign mem_0_89_W0_addr = W0_addr;
  assign mem_0_89_W0_clk = W0_clk;
  assign mem_0_89_W0_data = W0_data[719:712];
  assign mem_0_89_W0_en = W0_en;
  assign mem_0_89_W0_mask = W0_mask[89];
  assign mem_0_89_R0_addr = R0_addr;
  assign mem_0_89_R0_clk = R0_clk;
  assign mem_0_89_R0_en = R0_en;
  assign mem_0_90_W0_addr = W0_addr;
  assign mem_0_90_W0_clk = W0_clk;
  assign mem_0_90_W0_data = W0_data[727:720];
  assign mem_0_90_W0_en = W0_en;
  assign mem_0_90_W0_mask = W0_mask[90];
  assign mem_0_90_R0_addr = R0_addr;
  assign mem_0_90_R0_clk = R0_clk;
  assign mem_0_90_R0_en = R0_en;
  assign mem_0_91_W0_addr = W0_addr;
  assign mem_0_91_W0_clk = W0_clk;
  assign mem_0_91_W0_data = W0_data[735:728];
  assign mem_0_91_W0_en = W0_en;
  assign mem_0_91_W0_mask = W0_mask[91];
  assign mem_0_91_R0_addr = R0_addr;
  assign mem_0_91_R0_clk = R0_clk;
  assign mem_0_91_R0_en = R0_en;
  assign mem_0_92_W0_addr = W0_addr;
  assign mem_0_92_W0_clk = W0_clk;
  assign mem_0_92_W0_data = W0_data[743:736];
  assign mem_0_92_W0_en = W0_en;
  assign mem_0_92_W0_mask = W0_mask[92];
  assign mem_0_92_R0_addr = R0_addr;
  assign mem_0_92_R0_clk = R0_clk;
  assign mem_0_92_R0_en = R0_en;
  assign mem_0_93_W0_addr = W0_addr;
  assign mem_0_93_W0_clk = W0_clk;
  assign mem_0_93_W0_data = W0_data[751:744];
  assign mem_0_93_W0_en = W0_en;
  assign mem_0_93_W0_mask = W0_mask[93];
  assign mem_0_93_R0_addr = R0_addr;
  assign mem_0_93_R0_clk = R0_clk;
  assign mem_0_93_R0_en = R0_en;
  assign mem_0_94_W0_addr = W0_addr;
  assign mem_0_94_W0_clk = W0_clk;
  assign mem_0_94_W0_data = W0_data[759:752];
  assign mem_0_94_W0_en = W0_en;
  assign mem_0_94_W0_mask = W0_mask[94];
  assign mem_0_94_R0_addr = R0_addr;
  assign mem_0_94_R0_clk = R0_clk;
  assign mem_0_94_R0_en = R0_en;
  assign mem_0_95_W0_addr = W0_addr;
  assign mem_0_95_W0_clk = W0_clk;
  assign mem_0_95_W0_data = W0_data[767:760];
  assign mem_0_95_W0_en = W0_en;
  assign mem_0_95_W0_mask = W0_mask[95];
  assign mem_0_95_R0_addr = R0_addr;
  assign mem_0_95_R0_clk = R0_clk;
  assign mem_0_95_R0_en = R0_en;
  assign mem_0_96_W0_addr = W0_addr;
  assign mem_0_96_W0_clk = W0_clk;
  assign mem_0_96_W0_data = W0_data[775:768];
  assign mem_0_96_W0_en = W0_en;
  assign mem_0_96_W0_mask = W0_mask[96];
  assign mem_0_96_R0_addr = R0_addr;
  assign mem_0_96_R0_clk = R0_clk;
  assign mem_0_96_R0_en = R0_en;
  assign mem_0_97_W0_addr = W0_addr;
  assign mem_0_97_W0_clk = W0_clk;
  assign mem_0_97_W0_data = W0_data[783:776];
  assign mem_0_97_W0_en = W0_en;
  assign mem_0_97_W0_mask = W0_mask[97];
  assign mem_0_97_R0_addr = R0_addr;
  assign mem_0_97_R0_clk = R0_clk;
  assign mem_0_97_R0_en = R0_en;
  assign mem_0_98_W0_addr = W0_addr;
  assign mem_0_98_W0_clk = W0_clk;
  assign mem_0_98_W0_data = W0_data[791:784];
  assign mem_0_98_W0_en = W0_en;
  assign mem_0_98_W0_mask = W0_mask[98];
  assign mem_0_98_R0_addr = R0_addr;
  assign mem_0_98_R0_clk = R0_clk;
  assign mem_0_98_R0_en = R0_en;
  assign mem_0_99_W0_addr = W0_addr;
  assign mem_0_99_W0_clk = W0_clk;
  assign mem_0_99_W0_data = W0_data[799:792];
  assign mem_0_99_W0_en = W0_en;
  assign mem_0_99_W0_mask = W0_mask[99];
  assign mem_0_99_R0_addr = R0_addr;
  assign mem_0_99_R0_clk = R0_clk;
  assign mem_0_99_R0_en = R0_en;
  assign mem_0_100_W0_addr = W0_addr;
  assign mem_0_100_W0_clk = W0_clk;
  assign mem_0_100_W0_data = W0_data[807:800];
  assign mem_0_100_W0_en = W0_en;
  assign mem_0_100_W0_mask = W0_mask[100];
  assign mem_0_100_R0_addr = R0_addr;
  assign mem_0_100_R0_clk = R0_clk;
  assign mem_0_100_R0_en = R0_en;
  assign mem_0_101_W0_addr = W0_addr;
  assign mem_0_101_W0_clk = W0_clk;
  assign mem_0_101_W0_data = W0_data[815:808];
  assign mem_0_101_W0_en = W0_en;
  assign mem_0_101_W0_mask = W0_mask[101];
  assign mem_0_101_R0_addr = R0_addr;
  assign mem_0_101_R0_clk = R0_clk;
  assign mem_0_101_R0_en = R0_en;
  assign mem_0_102_W0_addr = W0_addr;
  assign mem_0_102_W0_clk = W0_clk;
  assign mem_0_102_W0_data = W0_data[823:816];
  assign mem_0_102_W0_en = W0_en;
  assign mem_0_102_W0_mask = W0_mask[102];
  assign mem_0_102_R0_addr = R0_addr;
  assign mem_0_102_R0_clk = R0_clk;
  assign mem_0_102_R0_en = R0_en;
  assign mem_0_103_W0_addr = W0_addr;
  assign mem_0_103_W0_clk = W0_clk;
  assign mem_0_103_W0_data = W0_data[831:824];
  assign mem_0_103_W0_en = W0_en;
  assign mem_0_103_W0_mask = W0_mask[103];
  assign mem_0_103_R0_addr = R0_addr;
  assign mem_0_103_R0_clk = R0_clk;
  assign mem_0_103_R0_en = R0_en;
  assign mem_0_104_W0_addr = W0_addr;
  assign mem_0_104_W0_clk = W0_clk;
  assign mem_0_104_W0_data = W0_data[839:832];
  assign mem_0_104_W0_en = W0_en;
  assign mem_0_104_W0_mask = W0_mask[104];
  assign mem_0_104_R0_addr = R0_addr;
  assign mem_0_104_R0_clk = R0_clk;
  assign mem_0_104_R0_en = R0_en;
  assign mem_0_105_W0_addr = W0_addr;
  assign mem_0_105_W0_clk = W0_clk;
  assign mem_0_105_W0_data = W0_data[847:840];
  assign mem_0_105_W0_en = W0_en;
  assign mem_0_105_W0_mask = W0_mask[105];
  assign mem_0_105_R0_addr = R0_addr;
  assign mem_0_105_R0_clk = R0_clk;
  assign mem_0_105_R0_en = R0_en;
  assign mem_0_106_W0_addr = W0_addr;
  assign mem_0_106_W0_clk = W0_clk;
  assign mem_0_106_W0_data = W0_data[855:848];
  assign mem_0_106_W0_en = W0_en;
  assign mem_0_106_W0_mask = W0_mask[106];
  assign mem_0_106_R0_addr = R0_addr;
  assign mem_0_106_R0_clk = R0_clk;
  assign mem_0_106_R0_en = R0_en;
  assign mem_0_107_W0_addr = W0_addr;
  assign mem_0_107_W0_clk = W0_clk;
  assign mem_0_107_W0_data = W0_data[863:856];
  assign mem_0_107_W0_en = W0_en;
  assign mem_0_107_W0_mask = W0_mask[107];
  assign mem_0_107_R0_addr = R0_addr;
  assign mem_0_107_R0_clk = R0_clk;
  assign mem_0_107_R0_en = R0_en;
  assign mem_0_108_W0_addr = W0_addr;
  assign mem_0_108_W0_clk = W0_clk;
  assign mem_0_108_W0_data = W0_data[871:864];
  assign mem_0_108_W0_en = W0_en;
  assign mem_0_108_W0_mask = W0_mask[108];
  assign mem_0_108_R0_addr = R0_addr;
  assign mem_0_108_R0_clk = R0_clk;
  assign mem_0_108_R0_en = R0_en;
  assign mem_0_109_W0_addr = W0_addr;
  assign mem_0_109_W0_clk = W0_clk;
  assign mem_0_109_W0_data = W0_data[879:872];
  assign mem_0_109_W0_en = W0_en;
  assign mem_0_109_W0_mask = W0_mask[109];
  assign mem_0_109_R0_addr = R0_addr;
  assign mem_0_109_R0_clk = R0_clk;
  assign mem_0_109_R0_en = R0_en;
  assign mem_0_110_W0_addr = W0_addr;
  assign mem_0_110_W0_clk = W0_clk;
  assign mem_0_110_W0_data = W0_data[887:880];
  assign mem_0_110_W0_en = W0_en;
  assign mem_0_110_W0_mask = W0_mask[110];
  assign mem_0_110_R0_addr = R0_addr;
  assign mem_0_110_R0_clk = R0_clk;
  assign mem_0_110_R0_en = R0_en;
  assign mem_0_111_W0_addr = W0_addr;
  assign mem_0_111_W0_clk = W0_clk;
  assign mem_0_111_W0_data = W0_data[895:888];
  assign mem_0_111_W0_en = W0_en;
  assign mem_0_111_W0_mask = W0_mask[111];
  assign mem_0_111_R0_addr = R0_addr;
  assign mem_0_111_R0_clk = R0_clk;
  assign mem_0_111_R0_en = R0_en;
  assign mem_0_112_W0_addr = W0_addr;
  assign mem_0_112_W0_clk = W0_clk;
  assign mem_0_112_W0_data = W0_data[903:896];
  assign mem_0_112_W0_en = W0_en;
  assign mem_0_112_W0_mask = W0_mask[112];
  assign mem_0_112_R0_addr = R0_addr;
  assign mem_0_112_R0_clk = R0_clk;
  assign mem_0_112_R0_en = R0_en;
  assign mem_0_113_W0_addr = W0_addr;
  assign mem_0_113_W0_clk = W0_clk;
  assign mem_0_113_W0_data = W0_data[911:904];
  assign mem_0_113_W0_en = W0_en;
  assign mem_0_113_W0_mask = W0_mask[113];
  assign mem_0_113_R0_addr = R0_addr;
  assign mem_0_113_R0_clk = R0_clk;
  assign mem_0_113_R0_en = R0_en;
  assign mem_0_114_W0_addr = W0_addr;
  assign mem_0_114_W0_clk = W0_clk;
  assign mem_0_114_W0_data = W0_data[919:912];
  assign mem_0_114_W0_en = W0_en;
  assign mem_0_114_W0_mask = W0_mask[114];
  assign mem_0_114_R0_addr = R0_addr;
  assign mem_0_114_R0_clk = R0_clk;
  assign mem_0_114_R0_en = R0_en;
  assign mem_0_115_W0_addr = W0_addr;
  assign mem_0_115_W0_clk = W0_clk;
  assign mem_0_115_W0_data = W0_data[927:920];
  assign mem_0_115_W0_en = W0_en;
  assign mem_0_115_W0_mask = W0_mask[115];
  assign mem_0_115_R0_addr = R0_addr;
  assign mem_0_115_R0_clk = R0_clk;
  assign mem_0_115_R0_en = R0_en;
  assign mem_0_116_W0_addr = W0_addr;
  assign mem_0_116_W0_clk = W0_clk;
  assign mem_0_116_W0_data = W0_data[935:928];
  assign mem_0_116_W0_en = W0_en;
  assign mem_0_116_W0_mask = W0_mask[116];
  assign mem_0_116_R0_addr = R0_addr;
  assign mem_0_116_R0_clk = R0_clk;
  assign mem_0_116_R0_en = R0_en;
  assign mem_0_117_W0_addr = W0_addr;
  assign mem_0_117_W0_clk = W0_clk;
  assign mem_0_117_W0_data = W0_data[943:936];
  assign mem_0_117_W0_en = W0_en;
  assign mem_0_117_W0_mask = W0_mask[117];
  assign mem_0_117_R0_addr = R0_addr;
  assign mem_0_117_R0_clk = R0_clk;
  assign mem_0_117_R0_en = R0_en;
  assign mem_0_118_W0_addr = W0_addr;
  assign mem_0_118_W0_clk = W0_clk;
  assign mem_0_118_W0_data = W0_data[951:944];
  assign mem_0_118_W0_en = W0_en;
  assign mem_0_118_W0_mask = W0_mask[118];
  assign mem_0_118_R0_addr = R0_addr;
  assign mem_0_118_R0_clk = R0_clk;
  assign mem_0_118_R0_en = R0_en;
  assign mem_0_119_W0_addr = W0_addr;
  assign mem_0_119_W0_clk = W0_clk;
  assign mem_0_119_W0_data = W0_data[959:952];
  assign mem_0_119_W0_en = W0_en;
  assign mem_0_119_W0_mask = W0_mask[119];
  assign mem_0_119_R0_addr = R0_addr;
  assign mem_0_119_R0_clk = R0_clk;
  assign mem_0_119_R0_en = R0_en;
  assign mem_0_120_W0_addr = W0_addr;
  assign mem_0_120_W0_clk = W0_clk;
  assign mem_0_120_W0_data = W0_data[967:960];
  assign mem_0_120_W0_en = W0_en;
  assign mem_0_120_W0_mask = W0_mask[120];
  assign mem_0_120_R0_addr = R0_addr;
  assign mem_0_120_R0_clk = R0_clk;
  assign mem_0_120_R0_en = R0_en;
  assign mem_0_121_W0_addr = W0_addr;
  assign mem_0_121_W0_clk = W0_clk;
  assign mem_0_121_W0_data = W0_data[975:968];
  assign mem_0_121_W0_en = W0_en;
  assign mem_0_121_W0_mask = W0_mask[121];
  assign mem_0_121_R0_addr = R0_addr;
  assign mem_0_121_R0_clk = R0_clk;
  assign mem_0_121_R0_en = R0_en;
  assign mem_0_122_W0_addr = W0_addr;
  assign mem_0_122_W0_clk = W0_clk;
  assign mem_0_122_W0_data = W0_data[983:976];
  assign mem_0_122_W0_en = W0_en;
  assign mem_0_122_W0_mask = W0_mask[122];
  assign mem_0_122_R0_addr = R0_addr;
  assign mem_0_122_R0_clk = R0_clk;
  assign mem_0_122_R0_en = R0_en;
  assign mem_0_123_W0_addr = W0_addr;
  assign mem_0_123_W0_clk = W0_clk;
  assign mem_0_123_W0_data = W0_data[991:984];
  assign mem_0_123_W0_en = W0_en;
  assign mem_0_123_W0_mask = W0_mask[123];
  assign mem_0_123_R0_addr = R0_addr;
  assign mem_0_123_R0_clk = R0_clk;
  assign mem_0_123_R0_en = R0_en;
  assign mem_0_124_W0_addr = W0_addr;
  assign mem_0_124_W0_clk = W0_clk;
  assign mem_0_124_W0_data = W0_data[999:992];
  assign mem_0_124_W0_en = W0_en;
  assign mem_0_124_W0_mask = W0_mask[124];
  assign mem_0_124_R0_addr = R0_addr;
  assign mem_0_124_R0_clk = R0_clk;
  assign mem_0_124_R0_en = R0_en;
  assign mem_0_125_W0_addr = W0_addr;
  assign mem_0_125_W0_clk = W0_clk;
  assign mem_0_125_W0_data = W0_data[1007:1000];
  assign mem_0_125_W0_en = W0_en;
  assign mem_0_125_W0_mask = W0_mask[125];
  assign mem_0_125_R0_addr = R0_addr;
  assign mem_0_125_R0_clk = R0_clk;
  assign mem_0_125_R0_en = R0_en;
  assign mem_0_126_W0_addr = W0_addr;
  assign mem_0_126_W0_clk = W0_clk;
  assign mem_0_126_W0_data = W0_data[1015:1008];
  assign mem_0_126_W0_en = W0_en;
  assign mem_0_126_W0_mask = W0_mask[126];
  assign mem_0_126_R0_addr = R0_addr;
  assign mem_0_126_R0_clk = R0_clk;
  assign mem_0_126_R0_en = R0_en;
  assign mem_0_127_W0_addr = W0_addr;
  assign mem_0_127_W0_clk = W0_clk;
  assign mem_0_127_W0_data = W0_data[1023:1016];
  assign mem_0_127_W0_en = W0_en;
  assign mem_0_127_W0_mask = W0_mask[127];
  assign mem_0_127_R0_addr = R0_addr;
  assign mem_0_127_R0_clk = R0_clk;
  assign mem_0_127_R0_en = R0_en;
  assign mem_0_128_W0_addr = W0_addr;
  assign mem_0_128_W0_clk = W0_clk;
  assign mem_0_128_W0_data = W0_data[1031:1024];
  assign mem_0_128_W0_en = W0_en;
  assign mem_0_128_W0_mask = W0_mask[128];
  assign mem_0_128_R0_addr = R0_addr;
  assign mem_0_128_R0_clk = R0_clk;
  assign mem_0_128_R0_en = R0_en;
  assign mem_0_129_W0_addr = W0_addr;
  assign mem_0_129_W0_clk = W0_clk;
  assign mem_0_129_W0_data = W0_data[1039:1032];
  assign mem_0_129_W0_en = W0_en;
  assign mem_0_129_W0_mask = W0_mask[129];
  assign mem_0_129_R0_addr = R0_addr;
  assign mem_0_129_R0_clk = R0_clk;
  assign mem_0_129_R0_en = R0_en;
  assign mem_0_130_W0_addr = W0_addr;
  assign mem_0_130_W0_clk = W0_clk;
  assign mem_0_130_W0_data = W0_data[1047:1040];
  assign mem_0_130_W0_en = W0_en;
  assign mem_0_130_W0_mask = W0_mask[130];
  assign mem_0_130_R0_addr = R0_addr;
  assign mem_0_130_R0_clk = R0_clk;
  assign mem_0_130_R0_en = R0_en;
  assign mem_0_131_W0_addr = W0_addr;
  assign mem_0_131_W0_clk = W0_clk;
  assign mem_0_131_W0_data = W0_data[1055:1048];
  assign mem_0_131_W0_en = W0_en;
  assign mem_0_131_W0_mask = W0_mask[131];
  assign mem_0_131_R0_addr = R0_addr;
  assign mem_0_131_R0_clk = R0_clk;
  assign mem_0_131_R0_en = R0_en;
  assign mem_0_132_W0_addr = W0_addr;
  assign mem_0_132_W0_clk = W0_clk;
  assign mem_0_132_W0_data = W0_data[1063:1056];
  assign mem_0_132_W0_en = W0_en;
  assign mem_0_132_W0_mask = W0_mask[132];
  assign mem_0_132_R0_addr = R0_addr;
  assign mem_0_132_R0_clk = R0_clk;
  assign mem_0_132_R0_en = R0_en;
  assign mem_0_133_W0_addr = W0_addr;
  assign mem_0_133_W0_clk = W0_clk;
  assign mem_0_133_W0_data = W0_data[1071:1064];
  assign mem_0_133_W0_en = W0_en;
  assign mem_0_133_W0_mask = W0_mask[133];
  assign mem_0_133_R0_addr = R0_addr;
  assign mem_0_133_R0_clk = R0_clk;
  assign mem_0_133_R0_en = R0_en;
  assign mem_0_134_W0_addr = W0_addr;
  assign mem_0_134_W0_clk = W0_clk;
  assign mem_0_134_W0_data = W0_data[1079:1072];
  assign mem_0_134_W0_en = W0_en;
  assign mem_0_134_W0_mask = W0_mask[134];
  assign mem_0_134_R0_addr = R0_addr;
  assign mem_0_134_R0_clk = R0_clk;
  assign mem_0_134_R0_en = R0_en;
  assign mem_0_135_W0_addr = W0_addr;
  assign mem_0_135_W0_clk = W0_clk;
  assign mem_0_135_W0_data = W0_data[1087:1080];
  assign mem_0_135_W0_en = W0_en;
  assign mem_0_135_W0_mask = W0_mask[135];
  assign mem_0_135_R0_addr = R0_addr;
  assign mem_0_135_R0_clk = R0_clk;
  assign mem_0_135_R0_en = R0_en;
  assign mem_0_136_W0_addr = W0_addr;
  assign mem_0_136_W0_clk = W0_clk;
  assign mem_0_136_W0_data = W0_data[1095:1088];
  assign mem_0_136_W0_en = W0_en;
  assign mem_0_136_W0_mask = W0_mask[136];
  assign mem_0_136_R0_addr = R0_addr;
  assign mem_0_136_R0_clk = R0_clk;
  assign mem_0_136_R0_en = R0_en;
  assign mem_0_137_W0_addr = W0_addr;
  assign mem_0_137_W0_clk = W0_clk;
  assign mem_0_137_W0_data = W0_data[1103:1096];
  assign mem_0_137_W0_en = W0_en;
  assign mem_0_137_W0_mask = W0_mask[137];
  assign mem_0_137_R0_addr = R0_addr;
  assign mem_0_137_R0_clk = R0_clk;
  assign mem_0_137_R0_en = R0_en;
  assign mem_0_138_W0_addr = W0_addr;
  assign mem_0_138_W0_clk = W0_clk;
  assign mem_0_138_W0_data = W0_data[1111:1104];
  assign mem_0_138_W0_en = W0_en;
  assign mem_0_138_W0_mask = W0_mask[138];
  assign mem_0_138_R0_addr = R0_addr;
  assign mem_0_138_R0_clk = R0_clk;
  assign mem_0_138_R0_en = R0_en;
  assign mem_0_139_W0_addr = W0_addr;
  assign mem_0_139_W0_clk = W0_clk;
  assign mem_0_139_W0_data = W0_data[1119:1112];
  assign mem_0_139_W0_en = W0_en;
  assign mem_0_139_W0_mask = W0_mask[139];
  assign mem_0_139_R0_addr = R0_addr;
  assign mem_0_139_R0_clk = R0_clk;
  assign mem_0_139_R0_en = R0_en;
  assign mem_0_140_W0_addr = W0_addr;
  assign mem_0_140_W0_clk = W0_clk;
  assign mem_0_140_W0_data = W0_data[1127:1120];
  assign mem_0_140_W0_en = W0_en;
  assign mem_0_140_W0_mask = W0_mask[140];
  assign mem_0_140_R0_addr = R0_addr;
  assign mem_0_140_R0_clk = R0_clk;
  assign mem_0_140_R0_en = R0_en;
  assign mem_0_141_W0_addr = W0_addr;
  assign mem_0_141_W0_clk = W0_clk;
  assign mem_0_141_W0_data = W0_data[1135:1128];
  assign mem_0_141_W0_en = W0_en;
  assign mem_0_141_W0_mask = W0_mask[141];
  assign mem_0_141_R0_addr = R0_addr;
  assign mem_0_141_R0_clk = R0_clk;
  assign mem_0_141_R0_en = R0_en;
  assign mem_0_142_W0_addr = W0_addr;
  assign mem_0_142_W0_clk = W0_clk;
  assign mem_0_142_W0_data = W0_data[1143:1136];
  assign mem_0_142_W0_en = W0_en;
  assign mem_0_142_W0_mask = W0_mask[142];
  assign mem_0_142_R0_addr = R0_addr;
  assign mem_0_142_R0_clk = R0_clk;
  assign mem_0_142_R0_en = R0_en;
  assign mem_0_143_W0_addr = W0_addr;
  assign mem_0_143_W0_clk = W0_clk;
  assign mem_0_143_W0_data = W0_data[1151:1144];
  assign mem_0_143_W0_en = W0_en;
  assign mem_0_143_W0_mask = W0_mask[143];
  assign mem_0_143_R0_addr = R0_addr;
  assign mem_0_143_R0_clk = R0_clk;
  assign mem_0_143_R0_en = R0_en;
  assign mem_0_144_W0_addr = W0_addr;
  assign mem_0_144_W0_clk = W0_clk;
  assign mem_0_144_W0_data = W0_data[1159:1152];
  assign mem_0_144_W0_en = W0_en;
  assign mem_0_144_W0_mask = W0_mask[144];
  assign mem_0_144_R0_addr = R0_addr;
  assign mem_0_144_R0_clk = R0_clk;
  assign mem_0_144_R0_en = R0_en;
  assign mem_0_145_W0_addr = W0_addr;
  assign mem_0_145_W0_clk = W0_clk;
  assign mem_0_145_W0_data = W0_data[1167:1160];
  assign mem_0_145_W0_en = W0_en;
  assign mem_0_145_W0_mask = W0_mask[145];
  assign mem_0_145_R0_addr = R0_addr;
  assign mem_0_145_R0_clk = R0_clk;
  assign mem_0_145_R0_en = R0_en;
  assign mem_0_146_W0_addr = W0_addr;
  assign mem_0_146_W0_clk = W0_clk;
  assign mem_0_146_W0_data = W0_data[1175:1168];
  assign mem_0_146_W0_en = W0_en;
  assign mem_0_146_W0_mask = W0_mask[146];
  assign mem_0_146_R0_addr = R0_addr;
  assign mem_0_146_R0_clk = R0_clk;
  assign mem_0_146_R0_en = R0_en;
  assign mem_0_147_W0_addr = W0_addr;
  assign mem_0_147_W0_clk = W0_clk;
  assign mem_0_147_W0_data = W0_data[1183:1176];
  assign mem_0_147_W0_en = W0_en;
  assign mem_0_147_W0_mask = W0_mask[147];
  assign mem_0_147_R0_addr = R0_addr;
  assign mem_0_147_R0_clk = R0_clk;
  assign mem_0_147_R0_en = R0_en;
  assign mem_0_148_W0_addr = W0_addr;
  assign mem_0_148_W0_clk = W0_clk;
  assign mem_0_148_W0_data = W0_data[1191:1184];
  assign mem_0_148_W0_en = W0_en;
  assign mem_0_148_W0_mask = W0_mask[148];
  assign mem_0_148_R0_addr = R0_addr;
  assign mem_0_148_R0_clk = R0_clk;
  assign mem_0_148_R0_en = R0_en;
  assign mem_0_149_W0_addr = W0_addr;
  assign mem_0_149_W0_clk = W0_clk;
  assign mem_0_149_W0_data = W0_data[1199:1192];
  assign mem_0_149_W0_en = W0_en;
  assign mem_0_149_W0_mask = W0_mask[149];
  assign mem_0_149_R0_addr = R0_addr;
  assign mem_0_149_R0_clk = R0_clk;
  assign mem_0_149_R0_en = R0_en;
  assign mem_0_150_W0_addr = W0_addr;
  assign mem_0_150_W0_clk = W0_clk;
  assign mem_0_150_W0_data = W0_data[1207:1200];
  assign mem_0_150_W0_en = W0_en;
  assign mem_0_150_W0_mask = W0_mask[150];
  assign mem_0_150_R0_addr = R0_addr;
  assign mem_0_150_R0_clk = R0_clk;
  assign mem_0_150_R0_en = R0_en;
  assign mem_0_151_W0_addr = W0_addr;
  assign mem_0_151_W0_clk = W0_clk;
  assign mem_0_151_W0_data = W0_data[1215:1208];
  assign mem_0_151_W0_en = W0_en;
  assign mem_0_151_W0_mask = W0_mask[151];
  assign mem_0_151_R0_addr = R0_addr;
  assign mem_0_151_R0_clk = R0_clk;
  assign mem_0_151_R0_en = R0_en;
  assign mem_0_152_W0_addr = W0_addr;
  assign mem_0_152_W0_clk = W0_clk;
  assign mem_0_152_W0_data = W0_data[1223:1216];
  assign mem_0_152_W0_en = W0_en;
  assign mem_0_152_W0_mask = W0_mask[152];
  assign mem_0_152_R0_addr = R0_addr;
  assign mem_0_152_R0_clk = R0_clk;
  assign mem_0_152_R0_en = R0_en;
  assign mem_0_153_W0_addr = W0_addr;
  assign mem_0_153_W0_clk = W0_clk;
  assign mem_0_153_W0_data = W0_data[1231:1224];
  assign mem_0_153_W0_en = W0_en;
  assign mem_0_153_W0_mask = W0_mask[153];
  assign mem_0_153_R0_addr = R0_addr;
  assign mem_0_153_R0_clk = R0_clk;
  assign mem_0_153_R0_en = R0_en;
  assign mem_0_154_W0_addr = W0_addr;
  assign mem_0_154_W0_clk = W0_clk;
  assign mem_0_154_W0_data = W0_data[1239:1232];
  assign mem_0_154_W0_en = W0_en;
  assign mem_0_154_W0_mask = W0_mask[154];
  assign mem_0_154_R0_addr = R0_addr;
  assign mem_0_154_R0_clk = R0_clk;
  assign mem_0_154_R0_en = R0_en;
  assign mem_0_155_W0_addr = W0_addr;
  assign mem_0_155_W0_clk = W0_clk;
  assign mem_0_155_W0_data = W0_data[1247:1240];
  assign mem_0_155_W0_en = W0_en;
  assign mem_0_155_W0_mask = W0_mask[155];
  assign mem_0_155_R0_addr = R0_addr;
  assign mem_0_155_R0_clk = R0_clk;
  assign mem_0_155_R0_en = R0_en;
  assign mem_0_156_W0_addr = W0_addr;
  assign mem_0_156_W0_clk = W0_clk;
  assign mem_0_156_W0_data = W0_data[1255:1248];
  assign mem_0_156_W0_en = W0_en;
  assign mem_0_156_W0_mask = W0_mask[156];
  assign mem_0_156_R0_addr = R0_addr;
  assign mem_0_156_R0_clk = R0_clk;
  assign mem_0_156_R0_en = R0_en;
  assign mem_0_157_W0_addr = W0_addr;
  assign mem_0_157_W0_clk = W0_clk;
  assign mem_0_157_W0_data = W0_data[1263:1256];
  assign mem_0_157_W0_en = W0_en;
  assign mem_0_157_W0_mask = W0_mask[157];
  assign mem_0_157_R0_addr = R0_addr;
  assign mem_0_157_R0_clk = R0_clk;
  assign mem_0_157_R0_en = R0_en;
  assign mem_0_158_W0_addr = W0_addr;
  assign mem_0_158_W0_clk = W0_clk;
  assign mem_0_158_W0_data = W0_data[1271:1264];
  assign mem_0_158_W0_en = W0_en;
  assign mem_0_158_W0_mask = W0_mask[158];
  assign mem_0_158_R0_addr = R0_addr;
  assign mem_0_158_R0_clk = R0_clk;
  assign mem_0_158_R0_en = R0_en;
  assign mem_0_159_W0_addr = W0_addr;
  assign mem_0_159_W0_clk = W0_clk;
  assign mem_0_159_W0_data = W0_data[1279:1272];
  assign mem_0_159_W0_en = W0_en;
  assign mem_0_159_W0_mask = W0_mask[159];
  assign mem_0_159_R0_addr = R0_addr;
  assign mem_0_159_R0_clk = R0_clk;
  assign mem_0_159_R0_en = R0_en;
  assign mem_0_160_W0_addr = W0_addr;
  assign mem_0_160_W0_clk = W0_clk;
  assign mem_0_160_W0_data = W0_data[1287:1280];
  assign mem_0_160_W0_en = W0_en;
  assign mem_0_160_W0_mask = W0_mask[160];
  assign mem_0_160_R0_addr = R0_addr;
  assign mem_0_160_R0_clk = R0_clk;
  assign mem_0_160_R0_en = R0_en;
  assign mem_0_161_W0_addr = W0_addr;
  assign mem_0_161_W0_clk = W0_clk;
  assign mem_0_161_W0_data = W0_data[1295:1288];
  assign mem_0_161_W0_en = W0_en;
  assign mem_0_161_W0_mask = W0_mask[161];
  assign mem_0_161_R0_addr = R0_addr;
  assign mem_0_161_R0_clk = R0_clk;
  assign mem_0_161_R0_en = R0_en;
  assign mem_0_162_W0_addr = W0_addr;
  assign mem_0_162_W0_clk = W0_clk;
  assign mem_0_162_W0_data = W0_data[1303:1296];
  assign mem_0_162_W0_en = W0_en;
  assign mem_0_162_W0_mask = W0_mask[162];
  assign mem_0_162_R0_addr = R0_addr;
  assign mem_0_162_R0_clk = R0_clk;
  assign mem_0_162_R0_en = R0_en;
  assign mem_0_163_W0_addr = W0_addr;
  assign mem_0_163_W0_clk = W0_clk;
  assign mem_0_163_W0_data = W0_data[1311:1304];
  assign mem_0_163_W0_en = W0_en;
  assign mem_0_163_W0_mask = W0_mask[163];
  assign mem_0_163_R0_addr = R0_addr;
  assign mem_0_163_R0_clk = R0_clk;
  assign mem_0_163_R0_en = R0_en;
  assign mem_0_164_W0_addr = W0_addr;
  assign mem_0_164_W0_clk = W0_clk;
  assign mem_0_164_W0_data = W0_data[1319:1312];
  assign mem_0_164_W0_en = W0_en;
  assign mem_0_164_W0_mask = W0_mask[164];
  assign mem_0_164_R0_addr = R0_addr;
  assign mem_0_164_R0_clk = R0_clk;
  assign mem_0_164_R0_en = R0_en;
  assign mem_0_165_W0_addr = W0_addr;
  assign mem_0_165_W0_clk = W0_clk;
  assign mem_0_165_W0_data = W0_data[1327:1320];
  assign mem_0_165_W0_en = W0_en;
  assign mem_0_165_W0_mask = W0_mask[165];
  assign mem_0_165_R0_addr = R0_addr;
  assign mem_0_165_R0_clk = R0_clk;
  assign mem_0_165_R0_en = R0_en;
  assign mem_0_166_W0_addr = W0_addr;
  assign mem_0_166_W0_clk = W0_clk;
  assign mem_0_166_W0_data = W0_data[1335:1328];
  assign mem_0_166_W0_en = W0_en;
  assign mem_0_166_W0_mask = W0_mask[166];
  assign mem_0_166_R0_addr = R0_addr;
  assign mem_0_166_R0_clk = R0_clk;
  assign mem_0_166_R0_en = R0_en;
  assign mem_0_167_W0_addr = W0_addr;
  assign mem_0_167_W0_clk = W0_clk;
  assign mem_0_167_W0_data = W0_data[1343:1336];
  assign mem_0_167_W0_en = W0_en;
  assign mem_0_167_W0_mask = W0_mask[167];
  assign mem_0_167_R0_addr = R0_addr;
  assign mem_0_167_R0_clk = R0_clk;
  assign mem_0_167_R0_en = R0_en;
  assign mem_0_168_W0_addr = W0_addr;
  assign mem_0_168_W0_clk = W0_clk;
  assign mem_0_168_W0_data = W0_data[1351:1344];
  assign mem_0_168_W0_en = W0_en;
  assign mem_0_168_W0_mask = W0_mask[168];
  assign mem_0_168_R0_addr = R0_addr;
  assign mem_0_168_R0_clk = R0_clk;
  assign mem_0_168_R0_en = R0_en;
  assign mem_0_169_W0_addr = W0_addr;
  assign mem_0_169_W0_clk = W0_clk;
  assign mem_0_169_W0_data = W0_data[1359:1352];
  assign mem_0_169_W0_en = W0_en;
  assign mem_0_169_W0_mask = W0_mask[169];
  assign mem_0_169_R0_addr = R0_addr;
  assign mem_0_169_R0_clk = R0_clk;
  assign mem_0_169_R0_en = R0_en;
  assign mem_0_170_W0_addr = W0_addr;
  assign mem_0_170_W0_clk = W0_clk;
  assign mem_0_170_W0_data = W0_data[1367:1360];
  assign mem_0_170_W0_en = W0_en;
  assign mem_0_170_W0_mask = W0_mask[170];
  assign mem_0_170_R0_addr = R0_addr;
  assign mem_0_170_R0_clk = R0_clk;
  assign mem_0_170_R0_en = R0_en;
  assign mem_0_171_W0_addr = W0_addr;
  assign mem_0_171_W0_clk = W0_clk;
  assign mem_0_171_W0_data = W0_data[1375:1368];
  assign mem_0_171_W0_en = W0_en;
  assign mem_0_171_W0_mask = W0_mask[171];
  assign mem_0_171_R0_addr = R0_addr;
  assign mem_0_171_R0_clk = R0_clk;
  assign mem_0_171_R0_en = R0_en;
  assign mem_0_172_W0_addr = W0_addr;
  assign mem_0_172_W0_clk = W0_clk;
  assign mem_0_172_W0_data = W0_data[1383:1376];
  assign mem_0_172_W0_en = W0_en;
  assign mem_0_172_W0_mask = W0_mask[172];
  assign mem_0_172_R0_addr = R0_addr;
  assign mem_0_172_R0_clk = R0_clk;
  assign mem_0_172_R0_en = R0_en;
  assign mem_0_173_W0_addr = W0_addr;
  assign mem_0_173_W0_clk = W0_clk;
  assign mem_0_173_W0_data = W0_data[1391:1384];
  assign mem_0_173_W0_en = W0_en;
  assign mem_0_173_W0_mask = W0_mask[173];
  assign mem_0_173_R0_addr = R0_addr;
  assign mem_0_173_R0_clk = R0_clk;
  assign mem_0_173_R0_en = R0_en;
  assign mem_0_174_W0_addr = W0_addr;
  assign mem_0_174_W0_clk = W0_clk;
  assign mem_0_174_W0_data = W0_data[1399:1392];
  assign mem_0_174_W0_en = W0_en;
  assign mem_0_174_W0_mask = W0_mask[174];
  assign mem_0_174_R0_addr = R0_addr;
  assign mem_0_174_R0_clk = R0_clk;
  assign mem_0_174_R0_en = R0_en;
  assign mem_0_175_W0_addr = W0_addr;
  assign mem_0_175_W0_clk = W0_clk;
  assign mem_0_175_W0_data = W0_data[1407:1400];
  assign mem_0_175_W0_en = W0_en;
  assign mem_0_175_W0_mask = W0_mask[175];
  assign mem_0_175_R0_addr = R0_addr;
  assign mem_0_175_R0_clk = R0_clk;
  assign mem_0_175_R0_en = R0_en;
  assign mem_0_176_W0_addr = W0_addr;
  assign mem_0_176_W0_clk = W0_clk;
  assign mem_0_176_W0_data = W0_data[1415:1408];
  assign mem_0_176_W0_en = W0_en;
  assign mem_0_176_W0_mask = W0_mask[176];
  assign mem_0_176_R0_addr = R0_addr;
  assign mem_0_176_R0_clk = R0_clk;
  assign mem_0_176_R0_en = R0_en;
  assign mem_0_177_W0_addr = W0_addr;
  assign mem_0_177_W0_clk = W0_clk;
  assign mem_0_177_W0_data = W0_data[1423:1416];
  assign mem_0_177_W0_en = W0_en;
  assign mem_0_177_W0_mask = W0_mask[177];
  assign mem_0_177_R0_addr = R0_addr;
  assign mem_0_177_R0_clk = R0_clk;
  assign mem_0_177_R0_en = R0_en;
  assign mem_0_178_W0_addr = W0_addr;
  assign mem_0_178_W0_clk = W0_clk;
  assign mem_0_178_W0_data = W0_data[1431:1424];
  assign mem_0_178_W0_en = W0_en;
  assign mem_0_178_W0_mask = W0_mask[178];
  assign mem_0_178_R0_addr = R0_addr;
  assign mem_0_178_R0_clk = R0_clk;
  assign mem_0_178_R0_en = R0_en;
  assign mem_0_179_W0_addr = W0_addr;
  assign mem_0_179_W0_clk = W0_clk;
  assign mem_0_179_W0_data = W0_data[1439:1432];
  assign mem_0_179_W0_en = W0_en;
  assign mem_0_179_W0_mask = W0_mask[179];
  assign mem_0_179_R0_addr = R0_addr;
  assign mem_0_179_R0_clk = R0_clk;
  assign mem_0_179_R0_en = R0_en;
  assign mem_0_180_W0_addr = W0_addr;
  assign mem_0_180_W0_clk = W0_clk;
  assign mem_0_180_W0_data = W0_data[1447:1440];
  assign mem_0_180_W0_en = W0_en;
  assign mem_0_180_W0_mask = W0_mask[180];
  assign mem_0_180_R0_addr = R0_addr;
  assign mem_0_180_R0_clk = R0_clk;
  assign mem_0_180_R0_en = R0_en;
  assign mem_0_181_W0_addr = W0_addr;
  assign mem_0_181_W0_clk = W0_clk;
  assign mem_0_181_W0_data = W0_data[1455:1448];
  assign mem_0_181_W0_en = W0_en;
  assign mem_0_181_W0_mask = W0_mask[181];
  assign mem_0_181_R0_addr = R0_addr;
  assign mem_0_181_R0_clk = R0_clk;
  assign mem_0_181_R0_en = R0_en;
  assign mem_0_182_W0_addr = W0_addr;
  assign mem_0_182_W0_clk = W0_clk;
  assign mem_0_182_W0_data = W0_data[1463:1456];
  assign mem_0_182_W0_en = W0_en;
  assign mem_0_182_W0_mask = W0_mask[182];
  assign mem_0_182_R0_addr = R0_addr;
  assign mem_0_182_R0_clk = R0_clk;
  assign mem_0_182_R0_en = R0_en;
  assign mem_0_183_W0_addr = W0_addr;
  assign mem_0_183_W0_clk = W0_clk;
  assign mem_0_183_W0_data = W0_data[1471:1464];
  assign mem_0_183_W0_en = W0_en;
  assign mem_0_183_W0_mask = W0_mask[183];
  assign mem_0_183_R0_addr = R0_addr;
  assign mem_0_183_R0_clk = R0_clk;
  assign mem_0_183_R0_en = R0_en;
  assign mem_0_184_W0_addr = W0_addr;
  assign mem_0_184_W0_clk = W0_clk;
  assign mem_0_184_W0_data = W0_data[1479:1472];
  assign mem_0_184_W0_en = W0_en;
  assign mem_0_184_W0_mask = W0_mask[184];
  assign mem_0_184_R0_addr = R0_addr;
  assign mem_0_184_R0_clk = R0_clk;
  assign mem_0_184_R0_en = R0_en;
  assign mem_0_185_W0_addr = W0_addr;
  assign mem_0_185_W0_clk = W0_clk;
  assign mem_0_185_W0_data = W0_data[1487:1480];
  assign mem_0_185_W0_en = W0_en;
  assign mem_0_185_W0_mask = W0_mask[185];
  assign mem_0_185_R0_addr = R0_addr;
  assign mem_0_185_R0_clk = R0_clk;
  assign mem_0_185_R0_en = R0_en;
  assign mem_0_186_W0_addr = W0_addr;
  assign mem_0_186_W0_clk = W0_clk;
  assign mem_0_186_W0_data = W0_data[1495:1488];
  assign mem_0_186_W0_en = W0_en;
  assign mem_0_186_W0_mask = W0_mask[186];
  assign mem_0_186_R0_addr = R0_addr;
  assign mem_0_186_R0_clk = R0_clk;
  assign mem_0_186_R0_en = R0_en;
  assign mem_0_187_W0_addr = W0_addr;
  assign mem_0_187_W0_clk = W0_clk;
  assign mem_0_187_W0_data = W0_data[1503:1496];
  assign mem_0_187_W0_en = W0_en;
  assign mem_0_187_W0_mask = W0_mask[187];
  assign mem_0_187_R0_addr = R0_addr;
  assign mem_0_187_R0_clk = R0_clk;
  assign mem_0_187_R0_en = R0_en;
  assign mem_0_188_W0_addr = W0_addr;
  assign mem_0_188_W0_clk = W0_clk;
  assign mem_0_188_W0_data = W0_data[1511:1504];
  assign mem_0_188_W0_en = W0_en;
  assign mem_0_188_W0_mask = W0_mask[188];
  assign mem_0_188_R0_addr = R0_addr;
  assign mem_0_188_R0_clk = R0_clk;
  assign mem_0_188_R0_en = R0_en;
  assign mem_0_189_W0_addr = W0_addr;
  assign mem_0_189_W0_clk = W0_clk;
  assign mem_0_189_W0_data = W0_data[1519:1512];
  assign mem_0_189_W0_en = W0_en;
  assign mem_0_189_W0_mask = W0_mask[189];
  assign mem_0_189_R0_addr = R0_addr;
  assign mem_0_189_R0_clk = R0_clk;
  assign mem_0_189_R0_en = R0_en;
  assign mem_0_190_W0_addr = W0_addr;
  assign mem_0_190_W0_clk = W0_clk;
  assign mem_0_190_W0_data = W0_data[1527:1520];
  assign mem_0_190_W0_en = W0_en;
  assign mem_0_190_W0_mask = W0_mask[190];
  assign mem_0_190_R0_addr = R0_addr;
  assign mem_0_190_R0_clk = R0_clk;
  assign mem_0_190_R0_en = R0_en;
  assign mem_0_191_W0_addr = W0_addr;
  assign mem_0_191_W0_clk = W0_clk;
  assign mem_0_191_W0_data = W0_data[1535:1528];
  assign mem_0_191_W0_en = W0_en;
  assign mem_0_191_W0_mask = W0_mask[191];
  assign mem_0_191_R0_addr = R0_addr;
  assign mem_0_191_R0_clk = R0_clk;
  assign mem_0_191_R0_en = R0_en;
  assign mem_0_192_W0_addr = W0_addr;
  assign mem_0_192_W0_clk = W0_clk;
  assign mem_0_192_W0_data = W0_data[1543:1536];
  assign mem_0_192_W0_en = W0_en;
  assign mem_0_192_W0_mask = W0_mask[192];
  assign mem_0_192_R0_addr = R0_addr;
  assign mem_0_192_R0_clk = R0_clk;
  assign mem_0_192_R0_en = R0_en;
  assign mem_0_193_W0_addr = W0_addr;
  assign mem_0_193_W0_clk = W0_clk;
  assign mem_0_193_W0_data = W0_data[1551:1544];
  assign mem_0_193_W0_en = W0_en;
  assign mem_0_193_W0_mask = W0_mask[193];
  assign mem_0_193_R0_addr = R0_addr;
  assign mem_0_193_R0_clk = R0_clk;
  assign mem_0_193_R0_en = R0_en;
  assign mem_0_194_W0_addr = W0_addr;
  assign mem_0_194_W0_clk = W0_clk;
  assign mem_0_194_W0_data = W0_data[1559:1552];
  assign mem_0_194_W0_en = W0_en;
  assign mem_0_194_W0_mask = W0_mask[194];
  assign mem_0_194_R0_addr = R0_addr;
  assign mem_0_194_R0_clk = R0_clk;
  assign mem_0_194_R0_en = R0_en;
  assign mem_0_195_W0_addr = W0_addr;
  assign mem_0_195_W0_clk = W0_clk;
  assign mem_0_195_W0_data = W0_data[1567:1560];
  assign mem_0_195_W0_en = W0_en;
  assign mem_0_195_W0_mask = W0_mask[195];
  assign mem_0_195_R0_addr = R0_addr;
  assign mem_0_195_R0_clk = R0_clk;
  assign mem_0_195_R0_en = R0_en;
  assign mem_0_196_W0_addr = W0_addr;
  assign mem_0_196_W0_clk = W0_clk;
  assign mem_0_196_W0_data = W0_data[1575:1568];
  assign mem_0_196_W0_en = W0_en;
  assign mem_0_196_W0_mask = W0_mask[196];
  assign mem_0_196_R0_addr = R0_addr;
  assign mem_0_196_R0_clk = R0_clk;
  assign mem_0_196_R0_en = R0_en;
  assign mem_0_197_W0_addr = W0_addr;
  assign mem_0_197_W0_clk = W0_clk;
  assign mem_0_197_W0_data = W0_data[1583:1576];
  assign mem_0_197_W0_en = W0_en;
  assign mem_0_197_W0_mask = W0_mask[197];
  assign mem_0_197_R0_addr = R0_addr;
  assign mem_0_197_R0_clk = R0_clk;
  assign mem_0_197_R0_en = R0_en;
  assign mem_0_198_W0_addr = W0_addr;
  assign mem_0_198_W0_clk = W0_clk;
  assign mem_0_198_W0_data = W0_data[1591:1584];
  assign mem_0_198_W0_en = W0_en;
  assign mem_0_198_W0_mask = W0_mask[198];
  assign mem_0_198_R0_addr = R0_addr;
  assign mem_0_198_R0_clk = R0_clk;
  assign mem_0_198_R0_en = R0_en;
  assign mem_0_199_W0_addr = W0_addr;
  assign mem_0_199_W0_clk = W0_clk;
  assign mem_0_199_W0_data = W0_data[1599:1592];
  assign mem_0_199_W0_en = W0_en;
  assign mem_0_199_W0_mask = W0_mask[199];
  assign mem_0_199_R0_addr = R0_addr;
  assign mem_0_199_R0_clk = R0_clk;
  assign mem_0_199_R0_en = R0_en;
  assign mem_0_200_W0_addr = W0_addr;
  assign mem_0_200_W0_clk = W0_clk;
  assign mem_0_200_W0_data = W0_data[1607:1600];
  assign mem_0_200_W0_en = W0_en;
  assign mem_0_200_W0_mask = W0_mask[200];
  assign mem_0_200_R0_addr = R0_addr;
  assign mem_0_200_R0_clk = R0_clk;
  assign mem_0_200_R0_en = R0_en;
  assign mem_0_201_W0_addr = W0_addr;
  assign mem_0_201_W0_clk = W0_clk;
  assign mem_0_201_W0_data = W0_data[1615:1608];
  assign mem_0_201_W0_en = W0_en;
  assign mem_0_201_W0_mask = W0_mask[201];
  assign mem_0_201_R0_addr = R0_addr;
  assign mem_0_201_R0_clk = R0_clk;
  assign mem_0_201_R0_en = R0_en;
  assign mem_0_202_W0_addr = W0_addr;
  assign mem_0_202_W0_clk = W0_clk;
  assign mem_0_202_W0_data = W0_data[1623:1616];
  assign mem_0_202_W0_en = W0_en;
  assign mem_0_202_W0_mask = W0_mask[202];
  assign mem_0_202_R0_addr = R0_addr;
  assign mem_0_202_R0_clk = R0_clk;
  assign mem_0_202_R0_en = R0_en;
  assign mem_0_203_W0_addr = W0_addr;
  assign mem_0_203_W0_clk = W0_clk;
  assign mem_0_203_W0_data = W0_data[1631:1624];
  assign mem_0_203_W0_en = W0_en;
  assign mem_0_203_W0_mask = W0_mask[203];
  assign mem_0_203_R0_addr = R0_addr;
  assign mem_0_203_R0_clk = R0_clk;
  assign mem_0_203_R0_en = R0_en;
  assign mem_0_204_W0_addr = W0_addr;
  assign mem_0_204_W0_clk = W0_clk;
  assign mem_0_204_W0_data = W0_data[1639:1632];
  assign mem_0_204_W0_en = W0_en;
  assign mem_0_204_W0_mask = W0_mask[204];
  assign mem_0_204_R0_addr = R0_addr;
  assign mem_0_204_R0_clk = R0_clk;
  assign mem_0_204_R0_en = R0_en;
  assign mem_0_205_W0_addr = W0_addr;
  assign mem_0_205_W0_clk = W0_clk;
  assign mem_0_205_W0_data = W0_data[1647:1640];
  assign mem_0_205_W0_en = W0_en;
  assign mem_0_205_W0_mask = W0_mask[205];
  assign mem_0_205_R0_addr = R0_addr;
  assign mem_0_205_R0_clk = R0_clk;
  assign mem_0_205_R0_en = R0_en;
  assign mem_0_206_W0_addr = W0_addr;
  assign mem_0_206_W0_clk = W0_clk;
  assign mem_0_206_W0_data = W0_data[1655:1648];
  assign mem_0_206_W0_en = W0_en;
  assign mem_0_206_W0_mask = W0_mask[206];
  assign mem_0_206_R0_addr = R0_addr;
  assign mem_0_206_R0_clk = R0_clk;
  assign mem_0_206_R0_en = R0_en;
  assign mem_0_207_W0_addr = W0_addr;
  assign mem_0_207_W0_clk = W0_clk;
  assign mem_0_207_W0_data = W0_data[1663:1656];
  assign mem_0_207_W0_en = W0_en;
  assign mem_0_207_W0_mask = W0_mask[207];
  assign mem_0_207_R0_addr = R0_addr;
  assign mem_0_207_R0_clk = R0_clk;
  assign mem_0_207_R0_en = R0_en;
  assign mem_0_208_W0_addr = W0_addr;
  assign mem_0_208_W0_clk = W0_clk;
  assign mem_0_208_W0_data = W0_data[1671:1664];
  assign mem_0_208_W0_en = W0_en;
  assign mem_0_208_W0_mask = W0_mask[208];
  assign mem_0_208_R0_addr = R0_addr;
  assign mem_0_208_R0_clk = R0_clk;
  assign mem_0_208_R0_en = R0_en;
  assign mem_0_209_W0_addr = W0_addr;
  assign mem_0_209_W0_clk = W0_clk;
  assign mem_0_209_W0_data = W0_data[1679:1672];
  assign mem_0_209_W0_en = W0_en;
  assign mem_0_209_W0_mask = W0_mask[209];
  assign mem_0_209_R0_addr = R0_addr;
  assign mem_0_209_R0_clk = R0_clk;
  assign mem_0_209_R0_en = R0_en;
  assign mem_0_210_W0_addr = W0_addr;
  assign mem_0_210_W0_clk = W0_clk;
  assign mem_0_210_W0_data = W0_data[1687:1680];
  assign mem_0_210_W0_en = W0_en;
  assign mem_0_210_W0_mask = W0_mask[210];
  assign mem_0_210_R0_addr = R0_addr;
  assign mem_0_210_R0_clk = R0_clk;
  assign mem_0_210_R0_en = R0_en;
  assign mem_0_211_W0_addr = W0_addr;
  assign mem_0_211_W0_clk = W0_clk;
  assign mem_0_211_W0_data = W0_data[1695:1688];
  assign mem_0_211_W0_en = W0_en;
  assign mem_0_211_W0_mask = W0_mask[211];
  assign mem_0_211_R0_addr = R0_addr;
  assign mem_0_211_R0_clk = R0_clk;
  assign mem_0_211_R0_en = R0_en;
  assign mem_0_212_W0_addr = W0_addr;
  assign mem_0_212_W0_clk = W0_clk;
  assign mem_0_212_W0_data = W0_data[1703:1696];
  assign mem_0_212_W0_en = W0_en;
  assign mem_0_212_W0_mask = W0_mask[212];
  assign mem_0_212_R0_addr = R0_addr;
  assign mem_0_212_R0_clk = R0_clk;
  assign mem_0_212_R0_en = R0_en;
  assign mem_0_213_W0_addr = W0_addr;
  assign mem_0_213_W0_clk = W0_clk;
  assign mem_0_213_W0_data = W0_data[1711:1704];
  assign mem_0_213_W0_en = W0_en;
  assign mem_0_213_W0_mask = W0_mask[213];
  assign mem_0_213_R0_addr = R0_addr;
  assign mem_0_213_R0_clk = R0_clk;
  assign mem_0_213_R0_en = R0_en;
  assign mem_0_214_W0_addr = W0_addr;
  assign mem_0_214_W0_clk = W0_clk;
  assign mem_0_214_W0_data = W0_data[1719:1712];
  assign mem_0_214_W0_en = W0_en;
  assign mem_0_214_W0_mask = W0_mask[214];
  assign mem_0_214_R0_addr = R0_addr;
  assign mem_0_214_R0_clk = R0_clk;
  assign mem_0_214_R0_en = R0_en;
  assign mem_0_215_W0_addr = W0_addr;
  assign mem_0_215_W0_clk = W0_clk;
  assign mem_0_215_W0_data = W0_data[1727:1720];
  assign mem_0_215_W0_en = W0_en;
  assign mem_0_215_W0_mask = W0_mask[215];
  assign mem_0_215_R0_addr = R0_addr;
  assign mem_0_215_R0_clk = R0_clk;
  assign mem_0_215_R0_en = R0_en;
  assign mem_0_216_W0_addr = W0_addr;
  assign mem_0_216_W0_clk = W0_clk;
  assign mem_0_216_W0_data = W0_data[1735:1728];
  assign mem_0_216_W0_en = W0_en;
  assign mem_0_216_W0_mask = W0_mask[216];
  assign mem_0_216_R0_addr = R0_addr;
  assign mem_0_216_R0_clk = R0_clk;
  assign mem_0_216_R0_en = R0_en;
  assign mem_0_217_W0_addr = W0_addr;
  assign mem_0_217_W0_clk = W0_clk;
  assign mem_0_217_W0_data = W0_data[1743:1736];
  assign mem_0_217_W0_en = W0_en;
  assign mem_0_217_W0_mask = W0_mask[217];
  assign mem_0_217_R0_addr = R0_addr;
  assign mem_0_217_R0_clk = R0_clk;
  assign mem_0_217_R0_en = R0_en;
  assign mem_0_218_W0_addr = W0_addr;
  assign mem_0_218_W0_clk = W0_clk;
  assign mem_0_218_W0_data = W0_data[1751:1744];
  assign mem_0_218_W0_en = W0_en;
  assign mem_0_218_W0_mask = W0_mask[218];
  assign mem_0_218_R0_addr = R0_addr;
  assign mem_0_218_R0_clk = R0_clk;
  assign mem_0_218_R0_en = R0_en;
  assign mem_0_219_W0_addr = W0_addr;
  assign mem_0_219_W0_clk = W0_clk;
  assign mem_0_219_W0_data = W0_data[1759:1752];
  assign mem_0_219_W0_en = W0_en;
  assign mem_0_219_W0_mask = W0_mask[219];
  assign mem_0_219_R0_addr = R0_addr;
  assign mem_0_219_R0_clk = R0_clk;
  assign mem_0_219_R0_en = R0_en;
  assign mem_0_220_W0_addr = W0_addr;
  assign mem_0_220_W0_clk = W0_clk;
  assign mem_0_220_W0_data = W0_data[1767:1760];
  assign mem_0_220_W0_en = W0_en;
  assign mem_0_220_W0_mask = W0_mask[220];
  assign mem_0_220_R0_addr = R0_addr;
  assign mem_0_220_R0_clk = R0_clk;
  assign mem_0_220_R0_en = R0_en;
  assign mem_0_221_W0_addr = W0_addr;
  assign mem_0_221_W0_clk = W0_clk;
  assign mem_0_221_W0_data = W0_data[1775:1768];
  assign mem_0_221_W0_en = W0_en;
  assign mem_0_221_W0_mask = W0_mask[221];
  assign mem_0_221_R0_addr = R0_addr;
  assign mem_0_221_R0_clk = R0_clk;
  assign mem_0_221_R0_en = R0_en;
  assign mem_0_222_W0_addr = W0_addr;
  assign mem_0_222_W0_clk = W0_clk;
  assign mem_0_222_W0_data = W0_data[1783:1776];
  assign mem_0_222_W0_en = W0_en;
  assign mem_0_222_W0_mask = W0_mask[222];
  assign mem_0_222_R0_addr = R0_addr;
  assign mem_0_222_R0_clk = R0_clk;
  assign mem_0_222_R0_en = R0_en;
  assign mem_0_223_W0_addr = W0_addr;
  assign mem_0_223_W0_clk = W0_clk;
  assign mem_0_223_W0_data = W0_data[1791:1784];
  assign mem_0_223_W0_en = W0_en;
  assign mem_0_223_W0_mask = W0_mask[223];
  assign mem_0_223_R0_addr = R0_addr;
  assign mem_0_223_R0_clk = R0_clk;
  assign mem_0_223_R0_en = R0_en;
  assign mem_0_224_W0_addr = W0_addr;
  assign mem_0_224_W0_clk = W0_clk;
  assign mem_0_224_W0_data = W0_data[1799:1792];
  assign mem_0_224_W0_en = W0_en;
  assign mem_0_224_W0_mask = W0_mask[224];
  assign mem_0_224_R0_addr = R0_addr;
  assign mem_0_224_R0_clk = R0_clk;
  assign mem_0_224_R0_en = R0_en;
  assign mem_0_225_W0_addr = W0_addr;
  assign mem_0_225_W0_clk = W0_clk;
  assign mem_0_225_W0_data = W0_data[1807:1800];
  assign mem_0_225_W0_en = W0_en;
  assign mem_0_225_W0_mask = W0_mask[225];
  assign mem_0_225_R0_addr = R0_addr;
  assign mem_0_225_R0_clk = R0_clk;
  assign mem_0_225_R0_en = R0_en;
  assign mem_0_226_W0_addr = W0_addr;
  assign mem_0_226_W0_clk = W0_clk;
  assign mem_0_226_W0_data = W0_data[1815:1808];
  assign mem_0_226_W0_en = W0_en;
  assign mem_0_226_W0_mask = W0_mask[226];
  assign mem_0_226_R0_addr = R0_addr;
  assign mem_0_226_R0_clk = R0_clk;
  assign mem_0_226_R0_en = R0_en;
  assign mem_0_227_W0_addr = W0_addr;
  assign mem_0_227_W0_clk = W0_clk;
  assign mem_0_227_W0_data = W0_data[1823:1816];
  assign mem_0_227_W0_en = W0_en;
  assign mem_0_227_W0_mask = W0_mask[227];
  assign mem_0_227_R0_addr = R0_addr;
  assign mem_0_227_R0_clk = R0_clk;
  assign mem_0_227_R0_en = R0_en;
  assign mem_0_228_W0_addr = W0_addr;
  assign mem_0_228_W0_clk = W0_clk;
  assign mem_0_228_W0_data = W0_data[1831:1824];
  assign mem_0_228_W0_en = W0_en;
  assign mem_0_228_W0_mask = W0_mask[228];
  assign mem_0_228_R0_addr = R0_addr;
  assign mem_0_228_R0_clk = R0_clk;
  assign mem_0_228_R0_en = R0_en;
  assign mem_0_229_W0_addr = W0_addr;
  assign mem_0_229_W0_clk = W0_clk;
  assign mem_0_229_W0_data = W0_data[1839:1832];
  assign mem_0_229_W0_en = W0_en;
  assign mem_0_229_W0_mask = W0_mask[229];
  assign mem_0_229_R0_addr = R0_addr;
  assign mem_0_229_R0_clk = R0_clk;
  assign mem_0_229_R0_en = R0_en;
  assign mem_0_230_W0_addr = W0_addr;
  assign mem_0_230_W0_clk = W0_clk;
  assign mem_0_230_W0_data = W0_data[1847:1840];
  assign mem_0_230_W0_en = W0_en;
  assign mem_0_230_W0_mask = W0_mask[230];
  assign mem_0_230_R0_addr = R0_addr;
  assign mem_0_230_R0_clk = R0_clk;
  assign mem_0_230_R0_en = R0_en;
  assign mem_0_231_W0_addr = W0_addr;
  assign mem_0_231_W0_clk = W0_clk;
  assign mem_0_231_W0_data = W0_data[1855:1848];
  assign mem_0_231_W0_en = W0_en;
  assign mem_0_231_W0_mask = W0_mask[231];
  assign mem_0_231_R0_addr = R0_addr;
  assign mem_0_231_R0_clk = R0_clk;
  assign mem_0_231_R0_en = R0_en;
  assign mem_0_232_W0_addr = W0_addr;
  assign mem_0_232_W0_clk = W0_clk;
  assign mem_0_232_W0_data = W0_data[1863:1856];
  assign mem_0_232_W0_en = W0_en;
  assign mem_0_232_W0_mask = W0_mask[232];
  assign mem_0_232_R0_addr = R0_addr;
  assign mem_0_232_R0_clk = R0_clk;
  assign mem_0_232_R0_en = R0_en;
  assign mem_0_233_W0_addr = W0_addr;
  assign mem_0_233_W0_clk = W0_clk;
  assign mem_0_233_W0_data = W0_data[1871:1864];
  assign mem_0_233_W0_en = W0_en;
  assign mem_0_233_W0_mask = W0_mask[233];
  assign mem_0_233_R0_addr = R0_addr;
  assign mem_0_233_R0_clk = R0_clk;
  assign mem_0_233_R0_en = R0_en;
  assign mem_0_234_W0_addr = W0_addr;
  assign mem_0_234_W0_clk = W0_clk;
  assign mem_0_234_W0_data = W0_data[1879:1872];
  assign mem_0_234_W0_en = W0_en;
  assign mem_0_234_W0_mask = W0_mask[234];
  assign mem_0_234_R0_addr = R0_addr;
  assign mem_0_234_R0_clk = R0_clk;
  assign mem_0_234_R0_en = R0_en;
  assign mem_0_235_W0_addr = W0_addr;
  assign mem_0_235_W0_clk = W0_clk;
  assign mem_0_235_W0_data = W0_data[1887:1880];
  assign mem_0_235_W0_en = W0_en;
  assign mem_0_235_W0_mask = W0_mask[235];
  assign mem_0_235_R0_addr = R0_addr;
  assign mem_0_235_R0_clk = R0_clk;
  assign mem_0_235_R0_en = R0_en;
  assign mem_0_236_W0_addr = W0_addr;
  assign mem_0_236_W0_clk = W0_clk;
  assign mem_0_236_W0_data = W0_data[1895:1888];
  assign mem_0_236_W0_en = W0_en;
  assign mem_0_236_W0_mask = W0_mask[236];
  assign mem_0_236_R0_addr = R0_addr;
  assign mem_0_236_R0_clk = R0_clk;
  assign mem_0_236_R0_en = R0_en;
  assign mem_0_237_W0_addr = W0_addr;
  assign mem_0_237_W0_clk = W0_clk;
  assign mem_0_237_W0_data = W0_data[1903:1896];
  assign mem_0_237_W0_en = W0_en;
  assign mem_0_237_W0_mask = W0_mask[237];
  assign mem_0_237_R0_addr = R0_addr;
  assign mem_0_237_R0_clk = R0_clk;
  assign mem_0_237_R0_en = R0_en;
  assign mem_0_238_W0_addr = W0_addr;
  assign mem_0_238_W0_clk = W0_clk;
  assign mem_0_238_W0_data = W0_data[1911:1904];
  assign mem_0_238_W0_en = W0_en;
  assign mem_0_238_W0_mask = W0_mask[238];
  assign mem_0_238_R0_addr = R0_addr;
  assign mem_0_238_R0_clk = R0_clk;
  assign mem_0_238_R0_en = R0_en;
  assign mem_0_239_W0_addr = W0_addr;
  assign mem_0_239_W0_clk = W0_clk;
  assign mem_0_239_W0_data = W0_data[1919:1912];
  assign mem_0_239_W0_en = W0_en;
  assign mem_0_239_W0_mask = W0_mask[239];
  assign mem_0_239_R0_addr = R0_addr;
  assign mem_0_239_R0_clk = R0_clk;
  assign mem_0_239_R0_en = R0_en;
  assign mem_0_240_W0_addr = W0_addr;
  assign mem_0_240_W0_clk = W0_clk;
  assign mem_0_240_W0_data = W0_data[1927:1920];
  assign mem_0_240_W0_en = W0_en;
  assign mem_0_240_W0_mask = W0_mask[240];
  assign mem_0_240_R0_addr = R0_addr;
  assign mem_0_240_R0_clk = R0_clk;
  assign mem_0_240_R0_en = R0_en;
  assign mem_0_241_W0_addr = W0_addr;
  assign mem_0_241_W0_clk = W0_clk;
  assign mem_0_241_W0_data = W0_data[1935:1928];
  assign mem_0_241_W0_en = W0_en;
  assign mem_0_241_W0_mask = W0_mask[241];
  assign mem_0_241_R0_addr = R0_addr;
  assign mem_0_241_R0_clk = R0_clk;
  assign mem_0_241_R0_en = R0_en;
  assign mem_0_242_W0_addr = W0_addr;
  assign mem_0_242_W0_clk = W0_clk;
  assign mem_0_242_W0_data = W0_data[1943:1936];
  assign mem_0_242_W0_en = W0_en;
  assign mem_0_242_W0_mask = W0_mask[242];
  assign mem_0_242_R0_addr = R0_addr;
  assign mem_0_242_R0_clk = R0_clk;
  assign mem_0_242_R0_en = R0_en;
  assign mem_0_243_W0_addr = W0_addr;
  assign mem_0_243_W0_clk = W0_clk;
  assign mem_0_243_W0_data = W0_data[1951:1944];
  assign mem_0_243_W0_en = W0_en;
  assign mem_0_243_W0_mask = W0_mask[243];
  assign mem_0_243_R0_addr = R0_addr;
  assign mem_0_243_R0_clk = R0_clk;
  assign mem_0_243_R0_en = R0_en;
  assign mem_0_244_W0_addr = W0_addr;
  assign mem_0_244_W0_clk = W0_clk;
  assign mem_0_244_W0_data = W0_data[1959:1952];
  assign mem_0_244_W0_en = W0_en;
  assign mem_0_244_W0_mask = W0_mask[244];
  assign mem_0_244_R0_addr = R0_addr;
  assign mem_0_244_R0_clk = R0_clk;
  assign mem_0_244_R0_en = R0_en;
  assign mem_0_245_W0_addr = W0_addr;
  assign mem_0_245_W0_clk = W0_clk;
  assign mem_0_245_W0_data = W0_data[1967:1960];
  assign mem_0_245_W0_en = W0_en;
  assign mem_0_245_W0_mask = W0_mask[245];
  assign mem_0_245_R0_addr = R0_addr;
  assign mem_0_245_R0_clk = R0_clk;
  assign mem_0_245_R0_en = R0_en;
  assign mem_0_246_W0_addr = W0_addr;
  assign mem_0_246_W0_clk = W0_clk;
  assign mem_0_246_W0_data = W0_data[1975:1968];
  assign mem_0_246_W0_en = W0_en;
  assign mem_0_246_W0_mask = W0_mask[246];
  assign mem_0_246_R0_addr = R0_addr;
  assign mem_0_246_R0_clk = R0_clk;
  assign mem_0_246_R0_en = R0_en;
  assign mem_0_247_W0_addr = W0_addr;
  assign mem_0_247_W0_clk = W0_clk;
  assign mem_0_247_W0_data = W0_data[1983:1976];
  assign mem_0_247_W0_en = W0_en;
  assign mem_0_247_W0_mask = W0_mask[247];
  assign mem_0_247_R0_addr = R0_addr;
  assign mem_0_247_R0_clk = R0_clk;
  assign mem_0_247_R0_en = R0_en;
  assign mem_0_248_W0_addr = W0_addr;
  assign mem_0_248_W0_clk = W0_clk;
  assign mem_0_248_W0_data = W0_data[1991:1984];
  assign mem_0_248_W0_en = W0_en;
  assign mem_0_248_W0_mask = W0_mask[248];
  assign mem_0_248_R0_addr = R0_addr;
  assign mem_0_248_R0_clk = R0_clk;
  assign mem_0_248_R0_en = R0_en;
  assign mem_0_249_W0_addr = W0_addr;
  assign mem_0_249_W0_clk = W0_clk;
  assign mem_0_249_W0_data = W0_data[1999:1992];
  assign mem_0_249_W0_en = W0_en;
  assign mem_0_249_W0_mask = W0_mask[249];
  assign mem_0_249_R0_addr = R0_addr;
  assign mem_0_249_R0_clk = R0_clk;
  assign mem_0_249_R0_en = R0_en;
  assign mem_0_250_W0_addr = W0_addr;
  assign mem_0_250_W0_clk = W0_clk;
  assign mem_0_250_W0_data = W0_data[2007:2000];
  assign mem_0_250_W0_en = W0_en;
  assign mem_0_250_W0_mask = W0_mask[250];
  assign mem_0_250_R0_addr = R0_addr;
  assign mem_0_250_R0_clk = R0_clk;
  assign mem_0_250_R0_en = R0_en;
  assign mem_0_251_W0_addr = W0_addr;
  assign mem_0_251_W0_clk = W0_clk;
  assign mem_0_251_W0_data = W0_data[2015:2008];
  assign mem_0_251_W0_en = W0_en;
  assign mem_0_251_W0_mask = W0_mask[251];
  assign mem_0_251_R0_addr = R0_addr;
  assign mem_0_251_R0_clk = R0_clk;
  assign mem_0_251_R0_en = R0_en;
  assign mem_0_252_W0_addr = W0_addr;
  assign mem_0_252_W0_clk = W0_clk;
  assign mem_0_252_W0_data = W0_data[2023:2016];
  assign mem_0_252_W0_en = W0_en;
  assign mem_0_252_W0_mask = W0_mask[252];
  assign mem_0_252_R0_addr = R0_addr;
  assign mem_0_252_R0_clk = R0_clk;
  assign mem_0_252_R0_en = R0_en;
  assign mem_0_253_W0_addr = W0_addr;
  assign mem_0_253_W0_clk = W0_clk;
  assign mem_0_253_W0_data = W0_data[2031:2024];
  assign mem_0_253_W0_en = W0_en;
  assign mem_0_253_W0_mask = W0_mask[253];
  assign mem_0_253_R0_addr = R0_addr;
  assign mem_0_253_R0_clk = R0_clk;
  assign mem_0_253_R0_en = R0_en;
  assign mem_0_254_W0_addr = W0_addr;
  assign mem_0_254_W0_clk = W0_clk;
  assign mem_0_254_W0_data = W0_data[2039:2032];
  assign mem_0_254_W0_en = W0_en;
  assign mem_0_254_W0_mask = W0_mask[254];
  assign mem_0_254_R0_addr = R0_addr;
  assign mem_0_254_R0_clk = R0_clk;
  assign mem_0_254_R0_en = R0_en;
  assign mem_0_255_W0_addr = W0_addr;
  assign mem_0_255_W0_clk = W0_clk;
  assign mem_0_255_W0_data = W0_data[2047:2040];
  assign mem_0_255_W0_en = W0_en;
  assign mem_0_255_W0_mask = W0_mask[255];
  assign mem_0_255_R0_addr = R0_addr;
  assign mem_0_255_R0_clk = R0_clk;
  assign mem_0_255_R0_en = R0_en;
endmodule
module tag_array_0_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [83:0] RW0_wdata,
  output [83:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [5:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [20:0] mem_0_0_RW0_wdata;
  wire [20:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [5:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [20:0] mem_0_1_RW0_wdata;
  wire [20:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [5:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [20:0] mem_0_2_RW0_wdata;
  wire [20:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [5:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [20:0] mem_0_3_RW0_wdata;
  wire [20:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [20:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [20:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [20:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [20:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [41:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [62:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [83:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [41:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [62:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_tag_array_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[20:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[41:21];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[62:42];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[83:63];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module data_arrays_0_0_ext(
  input  [7:0]   RW0_addr,
  input          RW0_clk,
  input  [127:0] RW0_wdata,
  output [127:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [3:0]   RW0_wmask
);
  wire [7:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [31:0] mem_0_0_RW0_wdata;
  wire [31:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [7:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [31:0] mem_0_1_RW0_wdata;
  wire [31:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [7:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [31:0] mem_0_2_RW0_wdata;
  wire [31:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [7:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [31:0] mem_0_3_RW0_wdata;
  wire [31:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [31:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [31:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [31:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [31:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [63:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [127:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [63:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_data_arrays_0_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[31:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[63:32];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[95:64];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[127:96];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module l2_tlb_ram_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [44:0] RW0_wdata,
  output [44:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [8:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [44:0] mem_0_0_RW0_wdata;
  wire [44:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire [44:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [44:0] RW0_rdata_0 = RW0_rdata_0_0;
  split_l2_tlb_ram_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata;
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata;
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
endmodule
module split_cc_dir_ext(
  input  [9:0]  RW0_addr,
  input         RW0_clk,
  input  [16:0] RW0_wdata,
  output [16:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] ram [0:1023];
  wire  ram_RW_0_r_en;
  wire [9:0] ram_RW_0_r_addr;
  wire [16:0] ram_RW_0_r_data;
  wire [16:0] ram_RW_0_w_data;
  wire [9:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[16:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_cc_banks_0_ext(
  input  [12:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:8191];
  wire  ram_RW_0_r_en;
  wire [12:0] ram_RW_0_r_addr;
  wire [63:0] ram_RW_0_r_data;
  wire [63:0] ram_RW_0_w_data;
  wire [12:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [12:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[12:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_data_arrays_0_ext(
  input  [7:0] RW0_addr,
  input        RW0_clk,
  input  [7:0] RW0_wdata,
  output [7:0] RW0_rdata,
  input        RW0_en,
  input        RW0_wmode,
  input        RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:255];
  wire  ram_RW_0_r_en;
  wire [7:0] ram_RW_0_r_addr;
  wire [7:0] ram_RW_0_r_data;
  wire [7:0] ram_RW_0_w_data;
  wire [7:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_tag_array_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [21:0] RW0_wdata,
  output [21:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] ram [0:63];
  wire  ram_RW_0_r_en;
  wire [5:0] ram_RW_0_r_addr;
  wire [21:0] ram_RW_0_r_data;
  wire [21:0] ram_RW_0_w_data;
  wire [5:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_mem_ext(
  input  [9:0] W0_addr,
  input        W0_clk,
  input  [7:0] W0_data,
  input        W0_en,
  input        W0_mask,
  input  [9:0] R0_addr,
  input        R0_clk,
  output [7:0] R0_data,
  input        R0_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:1023];
  wire  ram_R_0_en;
  wire [9:0] ram_R_0_addr;
  wire [7:0] ram_R_0_data;
  wire [7:0] ram_W_0_data;
  wire [9:0] ram_W_0_addr;
  wire  ram_W_0_mask;
  wire  ram_W_0_en;
  reg  ram_R_0_en_pipe_0;
  reg [9:0] ram_R_0_addr_pipe_0;
  assign ram_R_0_en = ram_R_0_en_pipe_0;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr];
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data;
  always @(posedge W0_clk) begin
    if (ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data;
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_mem_0_ext(
  input  [6:0] W0_addr,
  input        W0_clk,
  input  [7:0] W0_data,
  input        W0_en,
  input        W0_mask,
  input  [6:0] R0_addr,
  input        R0_clk,
  output [7:0] R0_data,
  input        R0_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127];
  wire  ram_R_0_en;
  wire [6:0] ram_R_0_addr;
  wire [7:0] ram_R_0_data;
  wire [7:0] ram_W_0_data;
  wire [6:0] ram_W_0_addr;
  wire  ram_W_0_mask;
  wire  ram_W_0_en;
  reg  ram_R_0_en_pipe_0;
  reg [6:0] ram_R_0_addr_pipe_0;
  assign ram_R_0_en = ram_R_0_en_pipe_0;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr];
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data;
  always @(posedge W0_clk) begin
    if (ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data;
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_tag_array_0_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [20:0] RW0_wdata,
  output [20:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] ram [0:63];
  wire  ram_RW_0_r_en;
  wire [5:0] ram_RW_0_r_addr;
  wire [20:0] ram_RW_0_r_data;
  wire [20:0] ram_RW_0_w_data;
  wire [5:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_data_arrays_0_0_ext(
  input  [7:0]  RW0_addr,
  input         RW0_clk,
  input  [31:0] RW0_wdata,
  output [31:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:255];
  wire  ram_RW_0_r_en;
  wire [7:0] ram_RW_0_r_addr;
  wire [31:0] ram_RW_0_r_data;
  wire [31:0] ram_RW_0_w_data;
  wire [7:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_l2_tlb_ram_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [44:0] RW0_wdata,
  output [44:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [44:0] ram [0:511];
  wire  ram_RW_0_r_en;
  wire [8:0] ram_RW_0_r_addr;
  wire [44:0] ram_RW_0_r_data;
  wire [44:0] ram_RW_0_w_data;
  wire [8:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [8:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[44:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
